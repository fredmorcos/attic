// FILE: FinalProcessor.vh

// ************************************************************************

// default verilog header file

// units of time and time resolution for this run
`timescale 1ps / 1ps

// this must be the very first module for interactive probing to work
module test;

// reg		a;
// wire		b;

// needed for interactive verilog probing.
   integer         tmp_channel;

// instantiate main verilog module
// NOTE: the name of the module must be the same as its type

	FinalProcessor FinalProcessor();

    initial
      begin
//    	$dumpfile();
//	$dumpvars;

//	a = 0;

// #1000 	a = 1; 

// #2000 	a = 0; 

//	$finish;
      end

endmodule

// include files
// `include "foo.v"

// ************************************************************************

// VERILOG netlist for "FinalProcessor" (generated by MMI_SUE4.4.0)

module DoubleInverter (in, out);
	input		in;
	output		out;
 
	wire		net_1;
 
	not #0 inv(net_1, in);
	not #0 inv_1(out, net_1);

endmodule		// DoubleInverter

module celltrans (in, out0, w);
	input		in;
	input		w;
	output		out0;
 
	wire		net_2;
	wire		net_1;
 
	not #0 inv(out0, net_2);
	not #0 inv_1(net_2, out0);
	not #0 inv_2(net_1, in);
	nmos n(net_2,net_1,w);

endmodule		// celltrans

module AluOrOutput (ALUOut, out);
	input	[31:0]	ALUOut;
	output		out;
 
	wire		net_28;
	wire		net_11;
	wire		net_30;
	wire		net_29;
	wire		net_12;
	wire		net_13;
	wire		net_14;
	wire		net_15;
	wire		net_16;
	wire		net_17;
	wire		net_18;
	wire		net_1;
	wire		net_20;
	wire		net_19;
	wire		net_2;
	wire		net_21;
	wire		net_3;
	wire		net_22;
	wire		net_4;
	wire		net_23;
	wire		net_5;
	wire		net_24;
	wire		net_6;
	wire		net_25;
	wire		net_7;
	wire		net_26;
	wire		net_8;
	wire		net_27;
	wire		net_10;
	wire		net_9;
 
	assign net_7 = !(ALUOut[12] || ALUOut[13]);
	assign net_30 = !(ALUOut[14] || ALUOut[15]);
	assign net_9 = !(net_7 || net_30);
	assign net_1 = !(ALUOut[8] || ALUOut[9]);
	assign net_12 = !(ALUOut[10] || ALUOut[11]);
	assign net_14 = !(net_1 || net_12);
	assign net_29 = !(ALUOut[4] || ALUOut[5]);
	assign net_16 = !(ALUOut[6] || ALUOut[7]);
	assign net_11 = !(net_29 || net_16);
	assign net_27 = !(ALUOut[0] || ALUOut[1]);
	assign net_24 = !(ALUOut[2] || ALUOut[3]);
	assign net_3 = !(net_27 || net_24);
	assign net_18 = !(ALUOut[28] || ALUOut[29]);
	assign net_6 = !(ALUOut[30] || ALUOut[31]);
	assign net_23 = !(net_18 || net_6);
	assign net_25 = !(ALUOut[24] || ALUOut[25]);
	assign net_28 = !(ALUOut[26] || ALUOut[27]);
	assign net_26 = !(net_25 || net_28);
	assign net_2 = !(ALUOut[20] || ALUOut[21]);
	assign net_20 = !(ALUOut[22] || ALUOut[23]);
	assign net_15 = !(net_2 || net_20);
	assign net_17 = !(ALUOut[16] || ALUOut[17]);
	assign net_8 = !(ALUOut[18] || ALUOut[19]);
	assign net_21 = !(net_17 || net_8);
	assign net_4 = !(net_26 || net_23);
	assign net_13 = !(net_21 || net_15);
	assign net_22 = !(net_14 || net_9);
	assign net_10 = !(net_3 || net_11);
	assign net_5 = !(net_13 || net_4);
	assign net_19 = !(net_10 || net_22);
	assign out = !(net_19 || net_5);

endmodule		// AluOrOutput

module Inverters32Bit (in, out);
	input	[31:0]	in;
	output	[31:0]	out;
 
	wire		net_28;
	wire		net_11;
	wire		net_30;
	wire		net_29;
	wire		net_12;
	wire		net_31;
	wire		net_13;
	wire		net_32;
	wire		net_14;
	wire		net_15;
	wire		net_16;
	wire		net_17;
	wire		net_18;
	wire		net_1;
	wire		net_20;
	wire		net_19;
	wire		net_2;
	wire		net_21;
	wire		net_3;
	wire		net_22;
	wire		net_4;
	wire		net_23;
	wire		net_5;
	wire		net_24;
	wire		net_6;
	wire		net_25;
	wire		net_7;
	wire		net_26;
	wire		net_8;
	wire		net_27;
	wire		net_10;
	wire		net_9;
 
	not #0 inv(net_13, in[0]);
	not #0 inv_1(out[0], net_13);
	not #0 inv_2(net_5, in[1]);
	not #0 inv_3(out[1], net_5);
	not #0 inv_4(net_18, in[2]);
	not #0 inv_5(out[2], net_18);
	not #0 inv_6(net_12, in[3]);
	not #0 inv_7(out[3], net_12);
	not #0 inv_8(net_4, in[4]);
	not #0 inv_9(out[4], net_4);
	not #0 inv_10(net_32, in[5]);
	not #0 inv_11(out[5], net_32);
	not #0 inv_12(net_29, in[6]);
	not #0 inv_13(out[6], net_29);
	not #0 inv_14(net_23, in[7]);
	not #0 inv_15(out[7], net_23);
	not #0 inv_16(net_8, in[8]);
	not #0 inv_17(out[8], net_8);
	not #0 inv_18(net_22, in[9]);
	not #0 inv_19(out[9], net_22);
	not #0 inv_20(net_11, in[10]);
	not #0 inv_21(out[10], net_11);
	not #0 inv_22(net_3, in[11]);
	not #0 inv_23(out[11], net_3);
	not #0 inv_24(net_9, in[12]);
	not #0 inv_25(out[12], net_9);
	not #0 inv_26(net_2, in[13]);
	not #0 inv_27(out[13], net_2);
	not #0 inv_28(net_31, in[14]);
	not #0 inv_29(out[14], net_31);
	not #0 inv_30(net_27, in[15]);
	not #0 inv_31(out[15], net_27);
	not #0 inv_32(net_20, in[16]);
	not #0 inv_33(out[16], net_20);
	not #0 inv_34(net_25, in[17]);
	not #0 inv_35(out[17], net_25);
	not #0 inv_36(net_16, in[18]);
	not #0 inv_37(out[18], net_16);
	not #0 inv_38(net_28, in[19]);
	not #0 inv_39(out[19], net_28);
	not #0 inv_40(net_21, in[20]);
	not #0 inv_41(out[20], net_21);
	not #0 inv_42(net_10, in[21]);
	not #0 inv_43(out[21], net_10);
	not #0 inv_44(net_19, in[22]);
	not #0 inv_45(out[22], net_19);
	not #0 inv_46(net_7, in[23]);
	not #0 inv_47(out[23], net_7);
	not #0 inv_48(net_24, in[24]);
	not #0 inv_49(out[24], net_24);
	not #0 inv_50(net_15, in[25]);
	not #0 inv_51(out[25], net_15);
	not #0 inv_52(net_1, in[26]);
	not #0 inv_53(out[26], net_1);
	not #0 inv_54(net_30, in[27]);
	not #0 inv_55(out[27], net_30);
	not #0 inv_56(net_26, in[28]);
	not #0 inv_57(out[28], net_26);
	not #0 inv_58(net_17, in[29]);
	not #0 inv_59(out[29], net_17);
	not #0 inv_60(net_6, in[30]);
	not #0 inv_61(out[30], net_6);
	not #0 inv_62(net_14, in[31]);
	not #0 inv_63(out[31], net_14);

endmodule		// Inverters32Bit

module pnzcell (alu, nout, pout, w, zout);
	input		w;
	input	[31:0]	alu;
	output		nout;
	output		pout;
	output		zout;
 
	wire		net_2;
	wire	[31:0]	ALU;
	wire		net_1;
 
	celltrans celltrans(.in(net_2), .out0(pout), .w(w));
	celltrans celltrans_1(.in(ALU[31]), .out0(nout), .w(w));
	celltrans celltrans_2(.in(net_1), .out0(zout), .w(w));
	AluOrOutput AluOrOutput(.out(net_1), .ALUOut(alu[31:0]));
	assign net_2 = !(ALU[31] || net_1);
	Inverters32Bit Inverters32Bit(.out(ALU[31:0]), .in(alu[31:0]));

endmodule		// pnzcell

module ripple8 (a, b, cin, cout, y);
	input		cin;
	input	[7:0]	a;
	input	[7:0]	b;
	output		cout;
	output	[7:0]	y;
 
	wire		net_1;
 
	ripple4 ripple4 (.b(b[7:4]), .a(a[7:4]), .cin(net_1), .sum(y[7:4]), 
		.cout(cout));
	ripple4 ripple4_1 (.b(b[3:0]), .a(a[3:0]), .cin(cin), .sum(y[3:0]), 
		.cout(net_1));

endmodule		// ripple8

module Adder32Bit (a, b, cin, cout, y);
	input		cin;
	input	[31:0]	a;
	input	[31:0]	b;
	output		cout;
	output	[31:0]	y;
 
	wire		net_2;
	wire		net_3;
	wire		net_1;
 
	ripple8 ripple8(.cout(net_1), .y(y[7:0]), .a(a[7:0]), .cin(cin), 
		.b(b[7:0]));
	ripple8 ripple8_1(.cin(net_2), .cout(net_3), .y(y[23:16]), 
		.a(a[23:16]), .b(b[23:16]));
	ripple8 ripple8_2(.cin(net_1), .cout(net_2), .y(y[15:8]), 
		.a(a[15:8]), .b(b[15:8]));
	ripple8 ripple8_3(.cin(net_3), .y(y[31:24]), .a(a[31:24]), 
		.b(b[31:24]), .cout(cout));

endmodule		// Adder32Bit

module Inverter32Bit (b, y);
	input	[31:0]	b;
	output	[31:0]	y;
 
	not #0 inv(y[0], b[0]);
	not #0 inv_1(y[1], b[1]);
	not #0 inv_2(y[2], b[2]);
	not #0 inv_3(y[3], b[3]);
	not #0 inv_4(y[4], b[4]);
	not #0 inv_5(y[5], b[5]);
	not #0 inv_6(y[6], b[6]);
	not #0 inv_7(y[7], b[7]);
	not #0 inv_8(y[8], b[8]);
	not #0 inv_9(y[9], b[9]);
	not #0 inv_10(y[10], b[10]);
	not #0 inv_11(y[11], b[11]);
	not #0 inv_12(y[12], b[12]);
	not #0 inv_13(y[13], b[13]);
	not #0 inv_14(y[14], b[14]);
	not #0 inv_15(y[15], b[15]);
	not #0 inv_16(y[16], b[16]);
	not #0 inv_17(y[17], b[17]);
	not #0 inv_18(y[18], b[18]);
	not #0 inv_19(y[19], b[19]);
	not #0 inv_20(y[20], b[20]);
	not #0 inv_21(y[21], b[21]);
	not #0 inv_22(y[22], b[22]);
	not #0 inv_23(y[23], b[23]);
	not #0 inv_24(y[24], b[24]);
	not #0 inv_25(y[25], b[25]);
	not #0 inv_26(y[26], b[26]);
	not #0 inv_27(y[27], b[27]);
	not #0 inv_28(y[28], b[28]);
	not #0 inv_29(y[29], b[29]);
	not #0 inv_30(y[30], b[30]);
	not #0 inv_31(y[31], b[31]);

endmodule		// Inverter32Bit

module Mux (a, b, s, y);
	input		a;
	input		b;
	input		s;
	output		y;
 
	wire		net_2;
	wire		net_3;
	wire		net_1;
 
	assign #0 net_3 = !(a && net_2);
	assign #0 net_1 = !(b && s);
	not #0 inv(net_2, s);
	assign #0 y = !(net_3 && net_1);

endmodule		// Mux

module Mux4Bit2to1 (a, b, s, y);
	input		s;
	input	[3:0]	a;
	input	[3:0]	b;
	output	[3:0]	y;
 
	wire		net_2;
	wire		net_1;
 
	Mux Mux(.s(net_2), .y(y[0]), .a(a[0]), .b(b[0]));
	Mux Mux_1(.s(net_2), .y(y[1]), .a(a[1]), .b(b[1]));
	Mux Mux_2(.s(net_2), .y(y[2]), .a(a[2]), .b(b[2]));
	Mux Mux_3(.s(net_2), .y(y[3]), .a(a[3]), .b(b[3]));
	not #0 inv(net_2, net_1);
	not #0 inv_1(net_1, s);

endmodule		// Mux4Bit2to1

module Mux32Bit2to1 (a, b, s, y);
	input		s;
	input	[31:0]	a;
	input	[31:0]	b;
	output	[31:0]	y;
 
	Mux4Bit2to1 Mux4Bit2to1(.y(y[3:0]), .a(a[3:0]), .b(b[3:0]), .s(s));
	Mux4Bit2to1 Mux4Bit2to1_1(.y(y[19:16]), .a(a[19:16]), .b(b[19:16]), 
		.s(s));
	Mux4Bit2to1 Mux4Bit2to1_2(.y(y[7:4]), .a(a[7:4]), .b(b[7:4]), .s(s));
	Mux4Bit2to1 Mux4Bit2to1_3(.y(y[23:20]), .a(a[23:20]), .b(b[23:20]), 
		.s(s));
	Mux4Bit2to1 Mux4Bit2to1_4(.y(y[11:8]), .a(a[11:8]), .b(b[11:8]), 
		.s(s));
	Mux4Bit2to1 Mux4Bit2to1_5(.y(y[27:24]), .a(a[27:24]), .b(b[27:24]), 
		.s(s));
	Mux4Bit2to1 Mux4Bit2to1_6(.y(y[15:12]), .a(a[15:12]), .b(b[15:12]), 
		.s(s));
	Mux4Bit2to1 Mux4Bit2to1_7(.y(y[31:28]), .a(a[31:28]), .b(b[31:28]), 
		.s(s));

endmodule		// Mux32Bit2to1

module Mux4to1 (a, b, c, d, s0, s1, y);
	input		a;
	input		b;
	input		c;
	input		d;
	input		s0;
	input		s1;
	output		y;
 
	wire		net_2;
	wire		net_1;
 
	Mux Mux(.y(net_2), .a(a), .b(b), .s(s0));
	Mux Mux_1(.y(net_1), .b(d), .s(s0), .a(c));
	Mux Mux_2(.b(net_1), .a(net_2), .s(s1), .y(y));

endmodule		// Mux4to1

module xgate (in, in_L, t1, t2);
	inout		t1;
	inout		t2;
	input		in;
	input		in_L;
 
	pmos p(t2,t1,in_L);
	nmos n(t2,t1,in);

endmodule		// xgate

module Hxor (in1, in2, out);
	input		in1;
	input		in2;
	output		out;
 
	wire		net_2;
	wire		net_3;
	wire		net_1;
 
	not #0 inv(net_3, in1);
	not #0 inv_1(out, net_2);
	not #0 inv_2(net_1, in2);
	xgate xgate(.t2(net_2), .in_L(net_3), .in(in1), .t1(in2));
	xgate xgate_1(.t1(net_1), .t2(net_2), .in(net_3), .in_L(in1));

endmodule		// Hxor

module Logic4Bit (a, b, s, y);
	input		a;
	input		b;
	input	[1:0]	s;
	output		y;
 
	wire		net_6;
	wire		net_2;
	wire		net_7;
	wire		net_3;
	wire		net_4;
	wire		net_5;
	wire		net_1;
 
	Mux4to1 Mux4to1(.d(net_1), .b(net_2), .c(net_3), .a(net_5), .y(y), 
		.s1(s[1]), .s0(s[0]));
	assign #0 net_7 = !(a && b);
	not #0 inv(net_5, net_7);
	assign net_6 = !(a || b);
	not #0 inv_1(net_2, net_6);
	not #0 inv_2(net_1, net_4);
	Hxor Hxor(.out(net_3), .in1(a), .in2(b));
	Hxor Hxor_1(.out(net_4), .in1(a), .in2(b));

endmodule		// Logic4Bit

module Logic32Bit (a, b, s, y);
	input	[31:0]	a;
	input	[31:0]	b;
	input	[1:0]	s;
	output	[31:0]	y;
 
	Logic4Bit Logic4Bit(.y(y[0]), .a(a[0]), .b(b[0]), .s(s[1:0]));
	Logic4Bit Logic4Bit_1(.y(y[1]), .a(a[1]), .b(b[1]), .s(s[1:0]));
	Logic4Bit Logic4Bit_2(.y(y[2]), .a(a[2]), .b(b[2]), .s(s[1:0]));
	Logic4Bit Logic4Bit_3(.y(y[3]), .a(a[3]), .b(b[3]), .s(s[1:0]));
	Logic4Bit Logic4Bit_4(.y(y[4]), .a(a[4]), .b(b[4]), .s(s[1:0]));
	Logic4Bit Logic4Bit_5(.y(y[5]), .a(a[5]), .b(b[5]), .s(s[1:0]));
	Logic4Bit Logic4Bit_6(.y(y[6]), .a(a[6]), .b(b[6]), .s(s[1:0]));
	Logic4Bit Logic4Bit_7(.y(y[7]), .a(a[7]), .b(b[7]), .s(s[1:0]));
	Logic4Bit Logic4Bit_8(.y(y[8]), .a(a[8]), .b(b[8]), .s(s[1:0]));
	Logic4Bit Logic4Bit_9(.y(y[9]), .a(a[9]), .b(b[9]), .s(s[1:0]));
	Logic4Bit Logic4Bit_10(.y(y[10]), .a(a[10]), .b(b[10]), .s(s[1:0]));
	Logic4Bit Logic4Bit_11(.y(y[11]), .a(a[11]), .b(b[11]), .s(s[1:0]));
	Logic4Bit Logic4Bit_12(.y(y[12]), .a(a[12]), .b(b[12]), .s(s[1:0]));
	Logic4Bit Logic4Bit_13(.y(y[13]), .a(a[13]), .b(b[13]), .s(s[1:0]));
	Logic4Bit Logic4Bit_14(.y(y[14]), .a(a[14]), .b(b[14]), .s(s[1:0]));
	Logic4Bit Logic4Bit_15(.y(y[15]), .a(a[15]), .b(b[15]), .s(s[1:0]));
	Logic4Bit Logic4Bit_16(.y(y[16]), .a(a[16]), .b(b[16]), .s(s[1:0]));
	Logic4Bit Logic4Bit_17(.y(y[17]), .a(a[17]), .b(b[17]), .s(s[1:0]));
	Logic4Bit Logic4Bit_18(.y(y[18]), .a(a[18]), .b(b[18]), .s(s[1:0]));
	Logic4Bit Logic4Bit_19(.y(y[19]), .a(a[19]), .b(b[19]), .s(s[1:0]));
	Logic4Bit Logic4Bit_20(.y(y[20]), .a(a[20]), .b(b[20]), .s(s[1:0]));
	Logic4Bit Logic4Bit_21(.y(y[21]), .a(a[21]), .b(b[21]), .s(s[1:0]));
	Logic4Bit Logic4Bit_22(.y(y[22]), .a(a[22]), .b(b[22]), .s(s[1:0]));
	Logic4Bit Logic4Bit_23(.y(y[23]), .a(a[23]), .b(b[23]), .s(s[1:0]));
	Logic4Bit Logic4Bit_24(.y(y[24]), .a(a[24]), .b(b[24]), .s(s[1:0]));
	Logic4Bit Logic4Bit_25(.y(y[25]), .a(a[25]), .b(b[25]), .s(s[1:0]));
	Logic4Bit Logic4Bit_26(.y(y[26]), .a(a[26]), .b(b[26]), .s(s[1:0]));
	Logic4Bit Logic4Bit_27(.y(y[27]), .a(a[27]), .b(b[27]), .s(s[1:0]));
	Logic4Bit Logic4Bit_28(.y(y[28]), .a(a[28]), .b(b[28]), .s(s[1:0]));
	Logic4Bit Logic4Bit_29(.y(y[29]), .a(a[29]), .b(b[29]), .s(s[1:0]));
	Logic4Bit Logic4Bit_30(.y(y[30]), .a(a[30]), .b(b[30]), .s(s[1:0]));
	Logic4Bit Logic4Bit_31(.y(y[31]), .a(a[31]), .b(b[31]), .s(s[1:0]));

endmodule		// Logic32Bit

module ALU (ALU_Result, a, b, overflow, s);
	input	[31:0]	a;
	input	[31:0]	b;
	input	[2:0]	s;
	output		overflow;
	output	[31:0]	ALU_Result;
 
	wire	[31:0]	net_2;
	wire	[31:0]	net_3;
	wire	[31:0]	net_4;
	wire	[31:0]	net_1;
 
	Adder32Bit Adder32Bit(.y(net_2[31:0]), .b(net_3[31:0]), 
		.cout(overflow), .a(a[31:0]), .cin(s[0]));
	Inverter32Bit Inverter32Bit(.y(net_1[31:0]), .b(b[31:0]));
	Mux32Bit2to1 Mux32Bit2to1(.b(net_1[31:0]), .y(net_3[31:0]), 
		.a(b[31:0]), .s(s[1]));
	Logic32Bit Logic32Bit(.y(net_4[31:0]), .a(a[31:0]), .b(b[31:0]), 
		.s(s[1:0]));
	Mux32Bit2to1 Mux32Bit2to1_1(.a(net_2[31:0]), .b(net_4[31:0]), 
		.y(ALU_Result[31:0]), .s(s[2]));

endmodule		// ALU

module cell32trans (in, out, w);
	input		w;
	input	[31:0]	in;
	output	[31:0]	out;
 
	celltrans celltrans(.out0(out[0]), .in(in[0]), .w(w));
	celltrans celltrans_1(.out0(out[1]), .in(in[1]), .w(w));
	celltrans celltrans_2(.out0(out[2]), .in(in[2]), .w(w));
	celltrans celltrans_3(.out0(out[3]), .in(in[3]), .w(w));
	celltrans celltrans_4(.out0(out[4]), .in(in[4]), .w(w));
	celltrans celltrans_5(.out0(out[5]), .in(in[5]), .w(w));
	celltrans celltrans_6(.out0(out[6]), .in(in[6]), .w(w));
	celltrans celltrans_7(.out0(out[7]), .in(in[7]), .w(w));
	celltrans celltrans_8(.out0(out[8]), .in(in[8]), .w(w));
	celltrans celltrans_9(.out0(out[9]), .in(in[9]), .w(w));
	celltrans celltrans_10(.out0(out[10]), .in(in[10]), .w(w));
	celltrans celltrans_11(.out0(out[11]), .in(in[11]), .w(w));
	celltrans celltrans_12(.out0(out[12]), .in(in[12]), .w(w));
	celltrans celltrans_13(.out0(out[13]), .in(in[13]), .w(w));
	celltrans celltrans_14(.out0(out[14]), .in(in[14]), .w(w));
	celltrans celltrans_15(.out0(out[15]), .in(in[15]), .w(w));
	celltrans celltrans_16(.out0(out[16]), .in(in[16]), .w(w));
	celltrans celltrans_17(.out0(out[17]), .in(in[17]), .w(w));
	celltrans celltrans_18(.out0(out[18]), .in(in[18]), .w(w));
	celltrans celltrans_19(.out0(out[19]), .in(in[19]), .w(w));
	celltrans celltrans_20(.out0(out[20]), .in(in[20]), .w(w));
	celltrans celltrans_21(.out0(out[21]), .in(in[21]), .w(w));
	celltrans celltrans_22(.out0(out[22]), .in(in[22]), .w(w));
	celltrans celltrans_23(.out0(out[23]), .in(in[23]), .w(w));
	celltrans celltrans_24(.out0(out[24]), .in(in[24]), .w(w));
	celltrans celltrans_25(.out0(out[25]), .in(in[25]), .w(w));
	celltrans celltrans_26(.out0(out[26]), .in(in[26]), .w(w));
	celltrans celltrans_27(.out0(out[27]), .in(in[27]), .w(w));
	celltrans celltrans_28(.out0(out[28]), .in(in[28]), .w(w));
	celltrans celltrans_29(.out0(out[29]), .in(in[29]), .w(w));
	celltrans celltrans_30(.out0(out[30]), .in(in[30]), .w(w));
	celltrans celltrans_31(.out0(out[31]), .in(in[31]), .w(w));

endmodule		// cell32trans

module ALU_UNIT (ALU_OP, ALU_OVERFLOW, ALU_RESULT, LATCH_WE, N_OUT, 
		PNZ_WE, P_OUT, R1, R2, Z_OUT);
	input		LATCH_WE;
	input		PNZ_WE;
	input	[2:0]	ALU_OP;
	input	[31:0]	R1;
	input	[31:0]	R2;
	output		ALU_OVERFLOW;
	output		N_OUT;
	output		P_OUT;
	output		Z_OUT;
	output	[31:0]	ALU_RESULT;
 
	wire	[31:0]	net_1;
	wire	[31:0]	net_2;
 
	pnzcell pnzcell(.zout(Z_OUT), .nout(N_OUT), .pout(P_OUT), 
		.alu(ALU_RESULT[31:0]), .w(PNZ_WE));
	ALU ALU(.a(net_1[31:0]), .b(net_2[31:0]), .s(ALU_OP[2:0]), 
		.ALU_Result(ALU_RESULT[31:0]), .overflow(ALU_OVERFLOW));
	cell32trans cell32trans(.out(net_1[31:0]), .in(R1[31:0]), 
		.w(LATCH_WE));
	cell32trans cell32trans_1(.out(net_2[31:0]), .in(R2[31:0]), 
		.w(LATCH_WE));

endmodule		// ALU_UNIT

module Inverters15Bit (in, out);
	input	[14:0]	in;
	output	[14:0]	out;
 
	wire		net_11;
	wire		net_12;
	wire		net_13;
	wire		net_14;
	wire		net_15;
	wire		net_1;
	wire		net_2;
	wire		net_3;
	wire		net_4;
	wire		net_5;
	wire		net_6;
	wire		net_7;
	wire		net_8;
	wire		net_10;
	wire		net_9;
 
	not #0 inv(net_14, in[0]);
	not #0 inv_1(out[0], net_14);
	not #0 inv_2(net_12, in[1]);
	not #0 inv_3(out[1], net_12);
	not #0 inv_4(net_2, in[2]);
	not #0 inv_5(out[2], net_2);
	not #0 inv_6(net_6, in[3]);
	not #0 inv_7(out[3], net_6);
	not #0 inv_8(net_15, in[4]);
	not #0 inv_9(out[4], net_15);
	not #0 inv_10(net_10, in[5]);
	not #0 inv_11(out[5], net_10);
	not #0 inv_12(net_8, in[6]);
	not #0 inv_13(out[6], net_8);
	not #0 inv_14(net_3, in[7]);
	not #0 inv_15(out[7], net_3);
	not #0 inv_16(net_13, in[8]);
	not #0 inv_17(out[8], net_13);
	not #0 inv_18(net_4, in[9]);
	not #0 inv_19(out[9], net_4);
	not #0 inv_20(net_7, in[10]);
	not #0 inv_21(out[10], net_7);
	not #0 inv_22(net_1, in[11]);
	not #0 inv_23(out[11], net_1);
	not #0 inv_24(net_11, in[12]);
	not #0 inv_25(out[12], net_11);
	not #0 inv_26(net_9, in[13]);
	not #0 inv_27(out[13], net_9);
	not #0 inv_28(net_5, in[14]);
	not #0 inv_29(out[14], net_5);
	not #0 inv_30(net_14, in[0]);
	not #0 inv_31(out[0], net_14);
	not #0 inv_32(net_12, in[1]);
	not #0 inv_33(out[1], net_12);
	not #0 inv_34(net_2, in[2]);
	not #0 inv_35(out[2], net_2);
	not #0 inv_36(net_6, in[3]);
	not #0 inv_37(out[3], net_6);
	not #0 inv_38(net_15, in[4]);
	not #0 inv_39(out[4], net_15);
	not #0 inv_40(net_10, in[5]);
	not #0 inv_41(out[5], net_10);
	not #0 inv_42(net_8, in[6]);
	not #0 inv_43(out[6], net_8);
	not #0 inv_44(net_3, in[7]);
	not #0 inv_45(out[7], net_3);
	not #0 inv_46(net_13, in[8]);
	not #0 inv_47(out[8], net_13);
	not #0 inv_48(net_4, in[9]);
	not #0 inv_49(out[9], net_4);
	not #0 inv_50(net_7, in[10]);
	not #0 inv_51(out[10], net_7);
	not #0 inv_52(net_1, in[11]);
	not #0 inv_53(out[11], net_1);
	not #0 inv_54(net_11, in[12]);
	not #0 inv_55(out[12], net_11);
	not #0 inv_56(net_9, in[13]);
	not #0 inv_57(out[13], net_9);
	not #0 inv_58(net_5, in[14]);
	not #0 inv_59(out[14], net_5);

endmodule		// Inverters15Bit

module Adder3217 (a, b, cout, y);
	input	[16:0]	a;
	input	[31:0]	b;
	output		cout;
	output	[31:0]	y;
 
	wire		net_2;
	wire		net_3;
	wire		net_1;
 
	ripple8 ripple8(.cout(net_2), .a(a[7:0]), .y(y[7:0]), .cin(1'b0), 
		.b(b[7:0]));
	ripple8 ripple8_1(.cin(net_1), .cout(net_3), .a(a[23:16]), 
		.y(y[23:16]), .b(b[23:16]));
	ripple8 ripple8_2(.cout(net_1), .cin(net_2), .a(a[15:8]), 
		.y(y[15:8]), .b(b[15:8]));
	ripple8 ripple8_3(.cin(net_3), .a(a[31:24]), .y(y[31:24]), 
		.b(b[31:24]), .cout(cout));
	DoubleInverter DoubleInverter(.in(a[16]), .out(a[16]));
	Inverters15Bit Inverters15Bit(.out(a[31:17]), 
		.in({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}));
		

endmodule		// Adder3217

module CUMuxSelect (L, S, T0, T3, s);
	input		L;
	input		S;
	input		T0;
	input		T3;
	output	[1:0]	s;
 
	wire		net_2;
	wire		net_3;
	wire		net_4;
	wire		net_1;
 
	assign net_4 = !(L || S);
	not #0 inv(net_2, net_4);
	assign #0 net_1 = !(net_2 && T3);
	not #0 inv_1(s[1], net_1);
	not #0 inv_2(net_3, T0);
	not #0 inv_3(s[0], net_3);

endmodule		// CUMuxSelect

module LoadStoreModule (LOAD, LS_ADDRESS, LS_OVERFLOW, OFFSET, 
		R_BASE_VALUE, S, STORE, T0, T3);
	input		LOAD;
	input		STORE;
	input		T0;
	input		T3;
	input	[16:0]	OFFSET;
	input	[31:0]	R_BASE_VALUE;
	output		LS_OVERFLOW;
	output	[31:0]	LS_ADDRESS;
	output	[1:0]	S;
 
	Adder3217 Adder3217(.y(LS_ADDRESS[31:0]), .b(R_BASE_VALUE[31:0]), 
		.cout(LS_OVERFLOW), .a(OFFSET[16:0]));
	CUMuxSelect CUMuxSelect(.L(LOAD), .T0(T0), .S(STORE), .s(S[1:0]), 
		.T3(T3));

endmodule		// LoadStoreModule

module mux32bit221 (a, b, s, y);
	input		s;
	input	[31:0]	a;
	input	[31:0]	b;
	output	[31:0]	y;
 
	Mux4Bit2to1 Mux4Bit2to1(.y(y[3:0]), .a(a[3:0]), .b(b[3:0]), .s(s));
	Mux4Bit2to1 Mux4Bit2to1_1(.y(y[19:16]), .a(a[19:16]), .b(b[19:16]), 
		.s(s));
	Mux4Bit2to1 Mux4Bit2to1_2(.y(y[7:4]), .a(a[7:4]), .b(b[7:4]), .s(s));
	Mux4Bit2to1 Mux4Bit2to1_3(.y(y[23:20]), .a(a[23:20]), .b(b[23:20]), 
		.s(s));
	Mux4Bit2to1 Mux4Bit2to1_4(.y(y[11:8]), .a(a[11:8]), .b(b[11:8]), 
		.s(s));
	Mux4Bit2to1 Mux4Bit2to1_5(.y(y[27:24]), .a(a[27:24]), .b(b[27:24]), 
		.s(s));
	Mux4Bit2to1 Mux4Bit2to1_6(.y(y[15:12]), .a(a[15:12]), .b(b[15:12]), 
		.s(s));
	Mux4Bit2to1 Mux4Bit2to1_7(.y(y[31:28]), .a(a[31:28]), .b(b[31:28]), 
		.s(s));

endmodule		// mux32bit221

module cell (in, out0, r1, w);
	input		in;
	input		r1;
	input		w;
	output		out0;
 
	wire		net_2;
	wire		net_3;
	wire		net_1;
 
	not #0 inv(net_2, net_1);
	not #0 inv_1(net_1, net_2);
	not #0 inv_2(net_3, in);
	nmos n(net_1,net_3,w);
	nmos n_1(out0,net_2,r1);

endmodule		// cell

module cell32 (in, out0, r, w);
	input		r;
	input		w;
	input	[31:0]	in;
	output	[31:0]	out0;
 
	cell cell(.out0(out0[18]), .r1(r), .in(in[18]), .w(w));
	cell cell_1(.out0(out0[17]), .r1(r), .in(in[17]), .w(w));
	cell cell_2(.out0(out0[19]), .r1(r), .in(in[19]), .w(w));
	cell cell_3(.out0(out0[20]), .r1(r), .in(in[20]), .w(w));
	cell cell_4(.out0(out0[21]), .r1(r), .in(in[21]), .w(w));
	cell cell_5(.out0(out0[22]), .r1(r), .in(in[22]), .w(w));
	cell cell_6(.out0(out0[23]), .r1(r), .in(in[23]), .w(w));
	cell cell_7(.out0(out0[31]), .r1(r), .in(in[31]), .w(w));
	cell cell_8(.out0(out0[30]), .r1(r), .in(in[30]), .w(w));
	cell cell_9(.out0(out0[29]), .r1(r), .in(in[29]), .w(w));
	cell cell_10(.out0(out0[28]), .r1(r), .in(in[28]), .w(w));
	cell cell_11(.out0(out0[27]), .r1(r), .in(in[27]), .w(w));
	cell cell_12(.out0(out0[26]), .r1(r), .in(in[26]), .w(w));
	cell cell_13(.out0(out0[25]), .r1(r), .in(in[25]), .w(w));
	cell cell_14(.out0(out0[24]), .r1(r), .in(in[24]), .w(w));
	cell cell_15(.out0(out0[16]), .r1(r), .in(in[16]), .w(w));
	cell cell_16(.out0(out0[8]), .r1(r), .in(in[8]), .w(w));
	cell cell_17(.out0(out0[9]), .r1(r), .in(in[9]), .w(w));
	cell cell_18(.out0(out0[10]), .r1(r), .in(in[10]), .w(w));
	cell cell_19(.out0(out0[11]), .r1(r), .in(in[11]), .w(w));
	cell cell_20(.out0(out0[12]), .r1(r), .in(in[12]), .w(w));
	cell cell_21(.out0(out0[13]), .r1(r), .in(in[13]), .w(w));
	cell cell_22(.out0(out0[14]), .r1(r), .in(in[14]), .w(w));
	cell cell_23(.out0(out0[15]), .r1(r), .in(in[15]), .w(w));
	cell cell_24(.out0(out0[7]), .r1(r), .in(in[7]), .w(w));
	cell cell_25(.out0(out0[6]), .r1(r), .in(in[6]), .w(w));
	cell cell_26(.out0(out0[5]), .r1(r), .in(in[5]), .w(w));
	cell cell_27(.out0(out0[4]), .r1(r), .in(in[4]), .w(w));
	cell cell_28(.out0(out0[3]), .r1(r), .in(in[3]), .w(w));
	cell cell_29(.out0(out0[2]), .r1(r), .in(in[2]), .w(w));
	cell cell_30(.out0(out0[1]), .r1(r), .in(in[1]), .w(w));
	cell cell_31(.out0(out0[0]), .r1(r), .in(in[0]), .w(w));

endmodule		// cell32

module halfadder (a, b, cout, s);
	input		a;
	input		b;
	output		cout;
	output		s;
 
	wire		net_1;
 
	assign #0 net_1 = !(a && b);
	not #0 inv(cout, net_1);
	Hxor Hxor(.in1(a), .in2(b), .out(s));

endmodule		// halfadder

module pcincrement (a, overflow, s);
	input	[31:0]	a;
	output		overflow;
	output	[31:0]	s;
 
	wire		net_28;
	wire		net_11;
	wire		net_30;
	wire		net_29;
	wire		net_12;
	wire		net_31;
	wire		net_13;
	wire		net_14;
	wire		net_15;
	wire		net_16;
	wire		net_17;
	wire		net_18;
	wire		net_1;
	wire		net_20;
	wire		net_19;
	wire		net_2;
	wire		net_21;
	wire		net_3;
	wire		net_22;
	wire		net_4;
	wire		net_23;
	wire		net_5;
	wire		net_24;
	wire		net_6;
	wire		net_25;
	wire		net_7;
	wire		net_26;
	wire		net_8;
	wire		net_27;
	wire		net_10;
	wire		net_9;
 
	halfadder halfadder(.cout(net_23), .a(a[2]), .s(s[2]), .b(1'b1));
	halfadder halfadder_1(.cout(net_12), .b(net_23), .a(a[3]), .s(s[3]));
	halfadder halfadder_2(.cout(net_10), .b(net_12), .a(a[4]), .s(s[4]));
	halfadder halfadder_3(.b(net_10), .cout(net_17), .a(a[5]), .s(s[5]));
	halfadder halfadder_4(.cout(net_4), .b(net_17), .a(a[6]), .s(s[6]));
	halfadder halfadder_5(.b(net_4), .cout(net_6), .a(a[7]), .s(s[7]));
	halfadder halfadder_6(.b(net_6), .cout(net_14), .a(a[8]), .s(s[8]));
	halfadder halfadder_7(.b(net_14), .cout(net_22), .a(a[9]), .s(s[9]));
	halfadder halfadder_8(.cout(net_16), .b(net_22), .a(a[10]), 
		.s(s[10]));
	halfadder halfadder_9(.cout(net_1), .b(net_16), .a(a[11]), 
		.s(s[11]));
	halfadder halfadder_10(.b(net_1), .cout(net_11), .a(a[12]), 
		.s(s[12]));
	halfadder halfadder_11(.b(net_11), .cout(net_29), .a(a[13]), 
		.s(s[13]));
	halfadder halfadder_12(.cout(net_18), .b(net_29), .a(a[14]), 
		.s(s[14]));
	halfadder halfadder_13(.cout(net_3), .b(net_18), .a(a[15]), 
		.s(s[15]));
	halfadder halfadder_14(.b(net_3), .cout(net_26), .a(a[16]), 
		.s(s[16]));
	halfadder halfadder_15(.cout(net_19), .b(net_26), .a(a[17]), 
		.s(s[17]));
	halfadder halfadder_16(.cout(net_9), .b(net_19), .a(a[18]), 
		.s(s[18]));
	halfadder halfadder_17(.cout(net_8), .b(net_9), .a(a[19]), 
		.s(s[19]));
	halfadder halfadder_18(.b(net_8), .cout(net_30), .a(a[20]), 
		.s(s[20]));
	halfadder halfadder_19(.cout(net_28), .b(net_30), .a(a[21]), 
		.s(s[21]));
	halfadder halfadder_20(.cout(net_25), .b(net_28), .a(a[22]), 
		.s(s[22]));
	halfadder halfadder_21(.cout(net_7), .b(net_25), .a(a[23]), 
		.s(s[23]));
	halfadder halfadder_22(.cout(net_2), .b(net_7), .a(a[24]), 
		.s(s[24]));
	halfadder halfadder_23(.b(net_2), .cout(net_15), .a(a[25]), 
		.s(s[25]));
	halfadder halfadder_24(.b(net_15), .cout(net_27), .a(a[26]), 
		.s(s[26]));
	halfadder halfadder_25(.cout(net_21), .b(net_27), .a(a[27]), 
		.s(s[27]));
	halfadder halfadder_26(.cout(net_5), .b(net_21), .a(a[28]), 
		.s(s[28]));
	halfadder halfadder_27(.b(net_5), .cout(net_13), .a(a[29]), 
		.s(s[29]));
	halfadder halfadder_28(.b(net_13), .cout(net_20), .a(a[30]), 
		.s(s[30]));
	halfadder halfadder_29(.b(net_20), .a(a[31]), .s(s[31]), 
		.cout(overflow));
	not #0 inv(net_24, a[0]);
	not #0 inv_1(s[0], net_24);
	not #0 inv_2(net_31, a[1]);
	not #0 inv_3(s[1], net_31);

endmodule		// pcincrement

module programcounter (BT, clock, out, overflow, s);
	input		clock;
	input		s;
	input	[31:0]	BT;
	output		overflow;
	output	[31:0]	out;
 
	wire	[31:0]	net_2;
	wire	[31:0]	net_1;
 
	mux32bit221 mux32bit221(.a(net_1[31:0]), .y(net_2[31:0]), 
		.b(BT[31:0]), .s(s));
	cell32 cell32(.in(net_2[31:0]), .w(clock), .out0(out[31:0]), 
		.r(1'b1));
	pcincrement pcincrement(.s(net_1[31:0]), .overflow(overflow), 
		.a(out[31:0]));

endmodule		// programcounter

module Flipflop (D, Q, clock_in, reset, reset_value);
	input		D;
	input		clock_in;
	input		reset;
	input		reset_value;
	output		Q;
 
	wire		net_6;
	wire		net_2;
	wire		net_3;
	wire		net_4;
	wire		net_5;
	wire		net_1;
 
	assign #0 net_3 = !(net_2 && net_1);
	assign #0 net_1 = !(net_3 && clock_in);
	assign #0 net_2 = !(net_4 && net_6);
	assign #0 Q = !(net_1 && net_5);
	assign #0 net_5 = !(Q && net_4);
	assign #0 net_4 = !(net_1 && clock_in && net_2);
	Mux Mux(.y(net_6), .a(D), .s(reset), .b(reset_value));

endmodule		// Flipflop

module SequenceCounter (CLOCK, T, reset);
	input		CLOCK;
	input		reset;
	output	[7:0]	T;
 
	Flipflop Flipflop(.clock_in(CLOCK), .Q(T[0]), .D(T[7]), 
		.reset(reset), .reset_value(1'b1));
	Flipflop Flipflop_1(.clock_in(CLOCK), .D(T[0]), .Q(T[1]), 
		.reset_value(1'b0), .reset(reset));
	Flipflop Flipflop_2(.clock_in(CLOCK), .D(T[1]), .Q(T[2]), 
		.reset_value(1'b0), .reset(reset));
	Flipflop Flipflop_3(.clock_in(CLOCK), .D(T[2]), .Q(T[3]), 
		.reset_value(1'b0), .reset(reset));
	Flipflop Flipflop_4(.clock_in(CLOCK), .D(T[3]), .Q(T[4]), 
		.reset_value(1'b0), .reset(reset));
	Flipflop Flipflop_5(.clock_in(CLOCK), .D(T[4]), .Q(T[5]), 
		.reset_value(1'b0), .reset(reset));
	Flipflop Flipflop_6(.clock_in(CLOCK), .D(T[5]), .Q(T[6]), 
		.reset_value(1'b0), .reset(reset));
	Flipflop Flipflop_7(.clock_in(CLOCK), .D(T[6]), .Q(T[7]), 
		.reset_value(1'b0), .reset(reset));

endmodule		// SequenceCounter

module decoder_2_4 (E, a, out);
	input		E;
	input	[1:0]	a;
	output	[3:0]	out;
 
	wire		net_6;
	wire		net_2;
	wire		net_7;
	wire		net_3;
	wire		net_8;
	wire		net_4;
	wire		net_5;
	wire		net_1;
 
	not #0 inv(net_5, a[0]);
	not #0 inv_1(net_4, a[1]);
	not #0 inv_2(net_7, a[0]);
	not #0 inv_3(net_6, a[1]);
	assign #0 net_2 = !(net_4 && net_5 && E);
	assign #0 net_1 = !(net_7 && a[1] && E);
	assign #0 net_3 = !(a[0] && net_6 && E);
	assign #0 net_8 = !(a[1] && a[0] && E);
	not #0 inv_4(out[0], net_2);
	not #0 inv_5(out[1], net_1);
	not #0 inv_6(out[2], net_3);
	not #0 inv_7(out[3], net_8);

endmodule		// decoder_2_4

module decoder_2_1_enable (a, e, out0, out1);
	input		a;
	input		e;
	output		out0;
	output		out1;
 
	wire		net_2;
	wire		net_3;
	wire		net_1;
 
	assign #0 net_3 = !(e && net_1);
	assign #0 net_2 = !(e && a);
	not #0 inv(out0, net_3);
	not #0 inv_1(out1, net_2);
	not #0 inv_2(net_1, a);

endmodule		// decoder_2_1_enable

module InstructionDecoder (ALU_UNIT_ACTIVATOR, BRANCH_UNIT_ACTIVATOR, 
		IR_OUT_27, IR_OUT_29, IR_OUT_30, IR_OUT_31, LOAD_UNIT_ACTIVATOR, 
		STORE_UNIT_ACTIVATOR);
	input		IR_OUT_27;
	input		IR_OUT_29;
	input		IR_OUT_30;
	input		IR_OUT_31;
	output		ALU_UNIT_ACTIVATOR;
	output		BRANCH_UNIT_ACTIVATOR;
	output		LOAD_UNIT_ACTIVATOR;
	output		STORE_UNIT_ACTIVATOR;
 
	wire	[3:0]	out;
	wire	[1:0]	t;
	wire		net_1;
	wire		net_2;
	wire		net_3;
	wire		net_4;
 
	Mux Mux(.y(t[0]), .b(IR_OUT_29), .a(IR_OUT_30), .s(IR_OUT_31));
	decoder_2_4 decoder_2_4(.out(out[3:0]), .a(t[1:0]), .E(vcc));
	decoder_2_1_enable decoder_2_1_enable(.e(out[2]), .a(IR_OUT_27), 
		.out1(STORE_UNIT_ACTIVATOR), .out0(LOAD_UNIT_ACTIVATOR));
	not #0 inv(t[1], net_4);
	not #0 inv_1(net_4, IR_OUT_31);
	not #0 inv_2(1'b0, net_3);
	not #0 inv_3(net_3, out[1]);
	not #0 inv_4(ALU_UNIT_ACTIVATOR, net_1);
	not #0 inv_5(net_1, out[0]);
	not #0 inv_6(BRANCH_UNIT_ACTIVATOR, net_2);
	not #0 inv_7(net_2, out[3]);

endmodule		// InstructionDecoder

module Inverters8Bits (in, out);
	input	[7:0]	in;
	output	[7:0]	out;
 
	wire		net_6;
	wire		net_2;
	wire		net_7;
	wire		net_3;
	wire		net_8;
	wire		net_4;
	wire		net_5;
	wire		net_1;
 
	not #0 inv(net_8, in[0]);
	not #0 inv_1(out[0], net_8);
	not #0 inv_2(net_1, in[1]);
	not #0 inv_3(out[1], net_1);
	not #0 inv_4(net_2, in[2]);
	not #0 inv_5(out[2], net_2);
	not #0 inv_6(net_4, in[3]);
	not #0 inv_7(out[3], net_4);
	not #0 inv_8(net_6, in[4]);
	not #0 inv_9(out[4], net_6);
	not #0 inv_10(net_3, in[5]);
	not #0 inv_11(out[5], net_3);
	not #0 inv_12(net_5, in[6]);
	not #0 inv_13(out[6], net_5);
	not #0 inv_14(net_7, in[7]);
	not #0 inv_15(out[7], net_7);

endmodule		// Inverters8Bits

module mux42132bbits (a, b, c, d, s, y);
	input	[31:0]	a;
	input	[31:0]	b;
	input	[31:0]	c;
	input	[31:0]	d;
	input	[1:0]	s;
	output	[31:0]	y;
 
	wire	[31:0]	net_2;
	wire	[31:0]	net_1;
 
	mux32bit221 mux32bit221(.y(net_1[31:0]), .a(a[31:0]), .b(b[31:0]), 
		.s(s[0]));
	mux32bit221 mux32bit221_1(.y(net_2[31:0]), .b(d[31:0]), .s(s[0]), 
		.a(c[31:0]));
	mux32bit221 mux32bit221_2(.a(net_1[31:0]), .b(net_2[31:0]), 
		.y(y[31:0]), .s(s[1]));

endmodule		// mux42132bbits

module controlunit (ADDRESS_SOURCE_SELECT, ALU_UNIT_ACTIVATOR, 
		BRANCH_ENABLE, BRANCH_TARGET, BRANCH_UNIT_ACTIVATOR, CLOCK, IR_OUT, 
		LOAD_UNIT_ACTIVATOR, LOAD_UNIT_ADDRESS, MAR_OUT, MAR_WE, MDR_IN, 
		MDR_OUT, MDR_WE, MDW_IN, MDW_OUT, MDW_WE, PC_OUT, PC_OVERFLOW, 
		SC_RESET, STORE_UNIT_ACTIVATOR, STORE_UNIT_ADDRESS, T_OUT);
	input		BRANCH_ENABLE;
	input		CLOCK;
	input		MAR_WE;
	input		MDR_WE;
	input		MDW_WE;
	input		SC_RESET;
	input	[1:0]	ADDRESS_SOURCE_SELECT;
	input	[31:0]	BRANCH_TARGET;
	input	[31:0]	LOAD_UNIT_ADDRESS;
	input	[31:0]	MDR_IN;
	input	[31:0]	MDW_IN;
	input	[31:0]	STORE_UNIT_ADDRESS;
	output		ALU_UNIT_ACTIVATOR;
	output		BRANCH_UNIT_ACTIVATOR;
	output		LOAD_UNIT_ACTIVATOR;
	output		PC_OVERFLOW;
	output		STORE_UNIT_ACTIVATOR;
	output	[31:0]	IR_OUT;
	output	[31:0]	MAR_OUT;
	output	[31:0]	MDR_OUT;
	output	[31:0]	MDW_OUT;
	output	[31:0]	PC_OUT;
	output	[7:0]	T_OUT;
 
	wire	[31:0]	IR;
	wire	[7:0]	T;
	wire	[31:0]	net_1;
	wire		net_2;
	wire		net_3;
 
	assign net_3 = !(T[0] || MAR_WE);
	not #0 inv(net_2, net_3);
	programcounter PC(.s(BRANCH_ENABLE), .clock(T[2]), 
		.overflow(PC_OVERFLOW), .out(PC_OUT[31:0]), 
		.BT(BRANCH_TARGET[31:0]));
	cell32trans cell32trans(.out(IR[31:0]), .w(T[2]), 
		.in(MDR_OUT[31:0]));
	cell32trans cell32trans_1(.in(MDR_IN[31:0]), .out(MDR_OUT[31:0]), 
		.w(MDR_WE));
	cell32trans cell32trans_2(.in(MDW_IN[31:0]), .w(MDW_WE), 
		.out(MDW_OUT[31:0]));
	cell32trans cell32trans_3(.in(net_1[31:0]), .w(net_2), 
		.out(MAR_OUT[31:0]));
	SequenceCounter SequenceCounter(.T(T[7:0]), .CLOCK(CLOCK), 
		.reset(SC_RESET));
	InstructionDecoder 
		InstructionDecoder(.BRANCH_UNIT_ACTIVATOR(BRANCH_UNIT_ACTIVATOR), 
		.IR_OUT_27(IR[27]), .IR_OUT_29(IR[29]), .IR_OUT_30(IR[30]), 
		.IR_OUT_31(IR[31]), .ALU_UNIT_ACTIVATOR(ALU_UNIT_ACTIVATOR), 
		.STORE_UNIT_ACTIVATOR(STORE_UNIT_ACTIVATOR), 
		.LOAD_UNIT_ACTIVATOR(LOAD_UNIT_ACTIVATOR));
	Inverters32Bit Inverters32Bit(.in(IR[31:0]), .out(IR_OUT[31:0]));
	Inverters8Bits Inverters8Bits(.in(T[7:0]), .out(T_OUT[7:0]));
	mux42132bbits mux42132bbits(.y(net_1[31:0]), 
		.s(ADDRESS_SOURCE_SELECT[1:0]), .c(STORE_UNIT_ADDRESS[31:0]), 
		.b(PC_OUT[31:0]), .d(LOAD_UNIT_ADDRESS[31:0]), .a(MAR_OUT[31:0]));

endmodule		// controlunit

module zero_register (out1, out2, r1, r2);
	input		r1;
	input		r2;
	output		out1;
	output		out2;
 
	nmos n(out1,1'b0,r1);
	nmos n_1(out2,1'b0,r2);

endmodule		// zero_register

module zero_32bit_register (out1, out2, r1, r2);
	input		r1;
	input		r2;
	output	[31:0]	out1;
	output	[31:0]	out2;
 
	zero_register zero_register(.r2(r2), .out1(out1[0]), .out2(out2[0]), 
		.r1(r1));
	zero_register zero_register_1(.r2(r2), .out1(out1[1]), 
		.out2(out2[1]), .r1(r1));
	zero_register zero_register_2(.r2(r2), .out1(out1[2]), 
		.out2(out2[2]), .r1(r1));
	zero_register zero_register_3(.r2(r2), .out1(out1[3]), 
		.out2(out2[3]), .r1(r1));
	zero_register zero_register_4(.r2(r2), .out1(out1[4]), 
		.out2(out2[4]), .r1(r1));
	zero_register zero_register_5(.r2(r2), .out1(out1[5]), 
		.out2(out2[5]), .r1(r1));
	zero_register zero_register_6(.r2(r2), .out1(out1[6]), 
		.out2(out2[6]), .r1(r1));
	zero_register zero_register_7(.r2(r2), .out1(out1[7]), 
		.out2(out2[7]), .r1(r1));
	zero_register zero_register_8(.r2(r2), .out1(out1[8]), 
		.out2(out2[8]), .r1(r1));
	zero_register zero_register_9(.r2(r2), .out1(out1[9]), 
		.out2(out2[9]), .r1(r1));
	zero_register zero_register_10(.r2(r2), .out1(out1[10]), 
		.out2(out2[10]), .r1(r1));
	zero_register zero_register_11(.r2(r2), .out1(out1[11]), 
		.out2(out2[11]), .r1(r1));
	zero_register zero_register_12(.r2(r2), .out1(out1[12]), 
		.out2(out2[12]), .r1(r1));
	zero_register zero_register_13(.r2(r2), .out1(out1[13]), 
		.out2(out2[13]), .r1(r1));
	zero_register zero_register_14(.r2(r2), .out1(out1[14]), 
		.out2(out2[14]), .r1(r1));
	zero_register zero_register_15(.r2(r2), .out1(out1[15]), 
		.out2(out2[15]), .r1(r1));
	zero_register zero_register_16(.r2(r2), .out1(out1[16]), 
		.out2(out2[16]), .r1(r1));
	zero_register zero_register_17(.r2(r2), .out1(out1[17]), 
		.out2(out2[17]), .r1(r1));
	zero_register zero_register_18(.r2(r2), .out1(out1[18]), 
		.out2(out2[18]), .r1(r1));
	zero_register zero_register_19(.r2(r2), .out1(out1[19]), 
		.out2(out2[19]), .r1(r1));
	zero_register zero_register_20(.r2(r2), .out1(out1[20]), 
		.out2(out2[20]), .r1(r1));
	zero_register zero_register_21(.r2(r2), .out1(out1[21]), 
		.out2(out2[21]), .r1(r1));
	zero_register zero_register_22(.r2(r2), .out1(out1[22]), 
		.out2(out2[22]), .r1(r1));
	zero_register zero_register_23(.r2(r2), .out1(out1[23]), 
		.out2(out2[23]), .r1(r1));
	zero_register zero_register_24(.r2(r2), .out1(out1[24]), 
		.out2(out2[24]), .r1(r1));
	zero_register zero_register_25(.r2(r2), .out1(out1[25]), 
		.out2(out2[25]), .r1(r1));
	zero_register zero_register_26(.r2(r2), .out1(out1[26]), 
		.out2(out2[26]), .r1(r1));
	zero_register zero_register_27(.r2(r2), .out1(out1[27]), 
		.out2(out2[27]), .r1(r1));
	zero_register zero_register_28(.r2(r2), .out1(out1[28]), 
		.out2(out2[28]), .r1(r1));
	zero_register zero_register_29(.r2(r2), .out1(out1[29]), 
		.out2(out2[29]), .r1(r1));
	zero_register zero_register_30(.r2(r2), .out1(out1[30]), 
		.out2(out2[30]), .r1(r1));
	zero_register zero_register_31(.r2(r2), .out1(out1[31]), 
		.out2(out2[31]), .r1(r1));

endmodule		// zero_32bit_register

module decoder_3_8 (out, s);
	input	[2:0]	s;
	output	[7:0]	out;
 
	wire		net_11;
	wire		net_12;
	wire		net_13;
	wire		net_14;
	wire		net_15;
	wire		net_16;
	wire		net_17;
	wire		net_18;
	wire		net_1;
	wire		net_20;
	wire		net_19;
	wire		net_2;
	wire		net_3;
	wire		net_4;
	wire		net_5;
	wire		net_6;
	wire		net_7;
	wire		net_8;
	wire		net_10;
	wire		net_9;
 
	not #0 inv(net_6, s[0]);
	not #0 inv_1(net_9, s[1]);
	not #0 inv_2(net_12, s[2]);
	not #0 inv_3(net_17, s[0]);
	not #0 inv_4(net_16, s[1]);
	not #0 inv_5(net_10, s[0]);
	not #0 inv_6(net_8, s[2]);
	not #0 inv_7(net_14, s[0]);
	not #0 inv_8(net_2, s[1]);
	not #0 inv_9(net_1, s[2]);
	not #0 inv_10(net_5, s[1]);
	not #0 inv_11(net_13, s[2]);
	not #0 inv_12(out[7], net_4);
	not #0 inv_13(out[6], net_19);
	not #0 inv_14(out[5], net_15);
	not #0 inv_15(out[4], net_7);
	not #0 inv_16(out[3], net_20);
	not #0 inv_17(out[2], net_18);
	not #0 inv_18(out[1], net_3);
	not #0 inv_19(out[0], net_11);
	assign #0 net_11 = !(net_6 && net_9 && net_12 && 1'b1);
	assign #0 net_4 = !(s[0] && s[1] && s[2] && 1'b1);
	assign #0 net_19 = !(s[0] && s[1] && net_13 && 1'b1);
	assign #0 net_15 = !(s[0] && net_5 && s[2] && 1'b1);
	assign #0 net_7 = !(s[0] && net_2 && net_1 && 1'b1);
	assign #0 net_20 = !(net_14 && s[1] && s[2] && 1'b1);
	assign #0 net_18 = !(net_10 && s[1] && net_8 && 1'b1);
	assign #0 net_3 = !(net_17 && net_16 && s[2] && 1'b1);

endmodule		// decoder_3_8

module decoder_5_32 (in, out);
	input	[4:0]	in;
	output	[31:0]	out;
 
	wire	[7:0]	dec_out;
 
	decoder_3_8 decoder_3_8(.out(dec_out[7:0]), .s(in[2:0]));
	decoder_2_4 decoder_2_4(.out(out[3:0]), .E(dec_out[0]), .a(in[4:3]));
	decoder_2_4 decoder_2_1(.out(out[7:4]), .E(dec_out[1]), .a(in[4:3]));
	decoder_2_4 decoder_2_2(.out(out[11:8]), .E(dec_out[2]), 
		.a(in[4:3]));
	decoder_2_4 decoder_2_3(.out(out[15:12]), .E(dec_out[3]), 
		.a(in[4:3]));
	decoder_2_4 decoder_2_5(.out(out[19:16]), .E(dec_out[4]), 
		.a(in[4:3]));
	decoder_2_4 decoder_2_6(.out(out[27:24]), .E(dec_out[6]), 
		.a(in[4:3]));
	decoder_2_4 decoder_2_7(.out(out[31:28]), .E(dec_out[7]), 
		.a(in[4:3]));
	decoder_2_4 decoder_2_8(.out(out[23:20]), .E(dec_out[5]), 
		.a(in[4:3]));

endmodule		// decoder_5_32

module write_enable (decoder_output, w, write_enable);
	input		write_enable;
	input	[31:1]	decoder_output;
	output	[31:1]	w;
 
	wire		net_28;
	wire		net_11;
	wire		net_30;
	wire		net_29;
	wire		net_12;
	wire		net_31;
	wire		net_13;
	wire		net_14;
	wire		net_15;
	wire		net_16;
	wire		net_17;
	wire		net_18;
	wire		net_1;
	wire		net_20;
	wire		net_19;
	wire		net_2;
	wire		net_21;
	wire		net_3;
	wire		net_22;
	wire		net_4;
	wire		net_23;
	wire		net_5;
	wire		net_24;
	wire		net_6;
	wire		net_25;
	wire		net_7;
	wire		net_26;
	wire		net_8;
	wire		net_27;
	wire		net_10;
	wire		net_9;
 
	assign #0 net_25 = !(decoder_output[1] && write_enable);
	not #0 inv(w[1], net_25);
	assign #0 net_18 = !(decoder_output[2] && write_enable);
	not #0 inv_1(w[2], net_18);
	assign #0 net_22 = !(decoder_output[3] && write_enable);
	not #0 inv_2(w[3], net_22);
	assign #0 net_27 = !(decoder_output[4] && write_enable);
	not #0 inv_3(w[4], net_27);
	assign #0 net_29 = !(decoder_output[5] && write_enable);
	not #0 inv_4(w[5], net_29);
	assign #0 net_31 = !(decoder_output[6] && write_enable);
	not #0 inv_5(w[6], net_31);
	assign #0 net_5 = !(decoder_output[7] && write_enable);
	not #0 inv_6(w[7], net_5);
	assign #0 net_1 = !(decoder_output[8] && write_enable);
	not #0 inv_7(w[8], net_1);
	assign #0 net_2 = !(decoder_output[9] && write_enable);
	not #0 inv_8(w[9], net_2);
	assign #0 net_6 = !(decoder_output[10] && write_enable);
	not #0 inv_9(w[10], net_6);
	assign #0 net_11 = !(decoder_output[11] && write_enable);
	not #0 inv_10(w[11], net_11);
	assign #0 net_13 = !(decoder_output[12] && write_enable);
	not #0 inv_11(w[12], net_13);
	assign #0 net_15 = !(decoder_output[13] && write_enable);
	not #0 inv_12(w[13], net_15);
	assign #0 net_16 = !(decoder_output[14] && write_enable);
	not #0 inv_13(w[14], net_16);
	assign #0 net_19 = !(decoder_output[15] && write_enable);
	not #0 inv_14(w[15], net_19);
	assign #0 net_23 = !(decoder_output[16] && write_enable);
	not #0 inv_15(w[16], net_23);
	assign #0 net_21 = !(decoder_output[17] && write_enable);
	not #0 inv_16(w[17], net_21);
	assign #0 net_24 = !(decoder_output[18] && write_enable);
	not #0 inv_17(w[18], net_24);
	assign #0 net_26 = !(decoder_output[19] && write_enable);
	not #0 inv_18(w[19], net_26);
	assign #0 net_28 = !(decoder_output[20] && write_enable);
	not #0 inv_19(w[20], net_28);
	assign #0 net_30 = !(decoder_output[21] && write_enable);
	not #0 inv_20(w[21], net_30);
	assign #0 net_4 = !(decoder_output[22] && write_enable);
	not #0 inv_21(w[22], net_4);
	assign #0 net_8 = !(decoder_output[23] && write_enable);
	not #0 inv_22(w[23], net_8);
	assign #0 net_10 = !(decoder_output[24] && write_enable);
	not #0 inv_23(w[24], net_10);
	assign #0 net_3 = !(decoder_output[25] && write_enable);
	not #0 inv_24(w[25], net_3);
	assign #0 net_7 = !(decoder_output[26] && write_enable);
	not #0 inv_25(w[26], net_7);
	assign #0 net_9 = !(decoder_output[27] && write_enable);
	not #0 inv_26(w[27], net_9);
	assign #0 net_12 = !(decoder_output[28] && write_enable);
	not #0 inv_27(w[28], net_12);
	assign #0 net_14 = !(decoder_output[29] && write_enable);
	not #0 inv_28(w[29], net_14);
	assign #0 net_17 = !(decoder_output[30] && write_enable);
	not #0 inv_29(w[30], net_17);
	assign #0 net_20 = !(decoder_output[31] && write_enable);
	not #0 inv_30(w[31], net_20);

endmodule		// write_enable

module register_32 (in, out1, out2, r1, r2, w);
	input		r1;
	input		r2;
	input		w;
	input	[31:0]	in;
	output	[31:0]	out1;
	output	[31:0]	out2;
 
	register_cell register_cell (.d(in[0]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[0]), .out2(out2[0]));
	register_cell register_cell_1 (.d(in[1]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[1]), .out2(out2[1]));
	register_cell register_cell_2 (.d(in[2]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[2]), .out2(out2[2]));
	register_cell register_cell_3 (.d(in[3]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[3]), .out2(out2[3]));
	register_cell register_cell_4 (.d(in[4]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[4]), .out2(out2[4]));
	register_cell register_cell_5 (.d(in[5]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[5]), .out2(out2[5]));
	register_cell register_cell_6 (.d(in[6]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[6]), .out2(out2[6]));
	register_cell register_cell_7 (.d(in[7]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[7]), .out2(out2[7]));
	register_cell register_cell_8 (.d(in[8]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[8]), .out2(out2[8]));
	register_cell register_cell_9 (.d(in[9]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[9]), .out2(out2[9]));
	register_cell register_cell_10 (.d(in[10]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[10]), .out2(out2[10]));
	register_cell register_cell_11 (.d(in[11]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[11]), .out2(out2[11]));
	register_cell register_cell_12 (.d(in[12]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[12]), .out2(out2[12]));
	register_cell register_cell_13 (.d(in[13]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[13]), .out2(out2[13]));
	register_cell register_cell_14 (.d(in[14]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[14]), .out2(out2[14]));
	register_cell register_cell_15 (.d(in[15]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[15]), .out2(out2[15]));
	register_cell register_cell_16 (.d(in[16]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[16]), .out2(out2[16]));
	register_cell register_cell_17 (.d(in[17]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[17]), .out2(out2[17]));
	register_cell register_cell_18 (.d(in[18]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[18]), .out2(out2[18]));
	register_cell register_cell_19 (.d(in[19]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[19]), .out2(out2[19]));
	register_cell register_cell_20 (.d(in[20]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[20]), .out2(out2[20]));
	register_cell register_cell_21 (.d(in[21]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[21]), .out2(out2[21]));
	register_cell register_cell_22 (.d(in[22]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[22]), .out2(out2[22]));
	register_cell register_cell_23 (.d(in[23]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[23]), .out2(out2[23]));
	register_cell register_cell_24 (.d(in[24]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[24]), .out2(out2[24]));
	register_cell register_cell_25 (.d(in[25]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[25]), .out2(out2[25]));
	register_cell register_cell_26 (.d(in[26]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[26]), .out2(out2[26]));
	register_cell register_cell_27 (.d(in[27]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[27]), .out2(out2[27]));
	register_cell register_cell_28 (.d(in[28]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[28]), .out2(out2[28]));
	register_cell register_cell_29 (.d(in[29]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[29]), .out2(out2[29]));
	register_cell register_cell_30 (.d(in[30]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[30]), .out2(out2[30]));
	register_cell register_cell_31 (.d(in[31]), .r1(r1), .r2(r2), .w(w), 
		.out1(out1[31]), .out2(out2[31]));

endmodule		// register_32

module Register_file_32bits (OUT1, OUT2, address_read1, address_read2, 
		address_write, data, write_enable);
	input		write_enable;
	input	[4:0]	address_read1;
	input	[4:0]	address_read2;
	input	[4:0]	address_write;
	input	[31:0]	data;
	output	[31:0]	OUT1;
	output	[31:0]	OUT2;
 
	wire	[31:0]	out1;
	wire	[31:0]	out2;
	wire	[31:0]	r1;
	wire	[31:0]	r2;
	wire	[13:13]	r3;
	wire	[31:1]	w;
	wire	[31:0]	dec_out;
 
	zero_32bit_register zero_32bit_register(.out1(out1[31:0]), 
		.out2(out2[31:0]), .r1(r1[0]), .r2(r2[0]));
	decoder_5_32 decoder_5_32(.out(r1[31:0]), .in(address_read1[4:0]));
	decoder_5_32 decoder_5_1(.out(r2[31:0]), .in(address_read2[4:0]));
	decoder_5_32 decoder_5_2(.in(address_write[4:0]), 
		.out(dec_out[31:0]));
	write_enable write_enable(.w(w[31:1]), .write_enable(write_enable), 
		.decoder_output(dec_out[31:1]));
	register_32 register_32(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[1]), .r2(r2[1]), .w(w[1]), .in(data[31:0]));
	register_32 register_1(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[2]), .r2(r2[2]), .w(w[2]), .in(data[31:0]));
	register_32 register_2(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[3]), .r2(r2[3]), .w(w[3]), .in(data[31:0]));
	register_32 register_3(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[4]), .r2(r2[4]), .w(w[4]), .in(data[31:0]));
	register_32 register_4(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[5]), .r2(r2[5]), .w(w[5]), .in(data[31:0]));
	register_32 register_5(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[6]), .r2(r2[6]), .w(w[6]), .in(data[31:0]));
	register_32 register_6(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[7]), .r2(r2[7]), .w(w[7]), .in(data[31:0]));
	register_32 register_7(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[8]), .r2(r2[8]), .w(w[8]), .in(data[31:0]));
	register_32 register_8(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[9]), .r2(r2[9]), .w(w[9]), .in(data[31:0]));
	register_32 register_9(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[10]), .r2(r2[10]), .w(w[10]), .in(data[31:0]));
	register_32 register_10(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[11]), .r2(r2[11]), .w(w[11]), .in(data[31:0]));
	register_32 register_11(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[12]), .r2(r2[12]), .w(w[12]), .in(data[31:0]));
	register_32 register_12(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[13]), .r2(r2[13]), .w(r3[13]), .in(data[31:0]));
	register_32 register_13(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[14]), .r2(r2[4]), .w(w[4]), .in(data[31:0]));
	register_32 register_14(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[15]), .r2(r2[15]), .w(w[15]), .in(data[31:0]));
	register_32 register_15(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[16]), .r2(r2[16]), .w(w[16]), .in(data[31:0]));
	register_32 register_16(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[17]), .r2(r2[17]), .w(w[17]), .in(data[31:0]));
	register_32 register_17(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[18]), .r2(r2[18]), .w(w[18]), .in(data[31:0]));
	register_32 register_18(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[19]), .r2(r2[19]), .w(w[19]), .in(data[31:0]));
	register_32 register_19(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[20]), .r2(r2[20]), .w(w[20]), .in(data[31:0]));
	register_32 register_20(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[21]), .r2(r2[21]), .w(w[21]), .in(data[31:0]));
	register_32 register_21(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[22]), .r2(r2[22]), .w(w[22]), .in(data[31:0]));
	register_32 register_22(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[23]), .r2(r2[23]), .w(w[23]), .in(data[31:0]));
	register_32 register_23(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[24]), .r2(r2[24]), .w(w[24]), .in(data[31:0]));
	register_32 register_24(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[25]), .r2(r2[25]), .w(w[25]), .in(data[31:0]));
	register_32 register_25(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[26]), .r2(r2[26]), .w(w[26]), .in(data[31:0]));
	register_32 register_26(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[27]), .r2(r2[27]), .w(w[27]), .in(data[31:0]));
	register_32 register_27(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[28]), .r2(r2[28]), .w(w[28]), .in(data[31:0]));
	register_32 register_28(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[29]), .r2(r2[29]), .w(w[29]), .in(data[31:0]));
	register_32 register_29(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[30]), .r2(r2[30]), .w(w[30]), .in(data[31:0]));
	register_32 register_30(.out1(out1[31:0]), .out2(out2[31:0]), 
		.r1(r1[31]), .r2(r2[31]), .w(w[31]), .in(data[31:0]));
	Inverters32Bit Inverters32Bit(.out(OUT1[31:0]), .in(out1[31:0]));
	Inverters32Bit Inverters32Bit_1(.out(OUT2[31:0]), .in(out2[31:0]));

endmodule		// Register_file_32bits

module FiveOnes (out);
	output	[4:0]	out;
 
	wire		net_2;
	wire		net_3;
	wire		net_4;
	wire		net_5;
	wire		net_1;
 
	not #0 inv(net_3, 1'b1);
	not #0 inv_1(out[0], net_3);
	not #0 inv_2(net_2, 1'b1);
	not #0 inv_3(out[1], net_2);
	not #0 inv_4(net_1, 1'b1);
	not #0 inv_5(out[2], net_1);
	not #0 inv_6(net_5, 1'b1);
	not #0 inv_7(out[3], net_5);
	not #0 inv_8(net_4, 1'b1);
	not #0 inv_9(out[4], net_4);

endmodule		// FiveOnes

module Mux32Bit8to1 (A, B, C, D, E, F, G, H, out, s);
	input	[31:0]	A;
	input	[31:0]	B;
	input	[31:0]	C;
	input	[31:0]	D;
	input	[31:0]	E;
	input	[31:0]	F;
	input	[31:0]	G;
	input	[31:0]	H;
	input	[2:0]	s;
	output	[31:0]	out;
 
	wire	[31:0]	net_1;
	wire	[31:0]	net_2;
 
	mux42132bbits mux42132bbits(.y(net_2[31:0]), .a(A[31:0]), 
		.b(B[31:0]), .s(s[1:0]), .c(C[31:0]), .d(D[31:0]));
	mux32bit221 mux32bit221(.b(net_1[31:0]), .a(net_2[31:0]), 
		.y(out[31:0]), .s(s[2]));
	mux42132bbits mux42132bbits_1(.y(net_1[31:0]), .s(s[1:0]), 
		.a(E[31:0]), .b(F[31:0]), .c(G[31:0]), .d(H[31:0]));

endmodule		// Mux32Bit8to1

module BranchDecoder (BC, BU, CallC, CallU, RetC, RetU, enable, s);
	input		enable;
	input	[2:0]	s;
	output		BC;
	output		BU;
	output		CallC;
	output		CallU;
	output		RetC;
	output		RetU;
 
	wire		net_11;
	wire		net_12;
	wire		net_13;
	wire		net_14;
	wire		net_15;
	wire		net_16;
	wire		net_17;
	wire		net_18;
	wire		net_1;
	wire		net_20;
	wire		net_19;
	wire		net_2;
	wire		net_3;
	wire		net_4;
	wire		net_5;
	wire		net_6;
	wire		net_7;
	wire		net_8;
	wire		net_10;
	wire		net_9;
 
	not #0 inv(net_4, s[0]);
	not #0 inv_1(net_17, s[1]);
	not #0 inv_2(net_9, s[2]);
	not #0 inv_3(net_15, s[0]);
	not #0 inv_4(net_7, s[1]);
	not #0 inv_5(net_1, s[0]);
	not #0 inv_6(net_3, s[2]);
	not #0 inv_7(net_13, s[0]);
	not #0 inv_8(net_5, s[1]);
	not #0 inv_9(net_8, s[2]);
	not #0 inv_10(net_14, s[1]);
	not #0 inv_11(net_10, s[2]);
	not #0 inv_12(1'b0, net_6);
	not #0 inv_13(1'b0, net_20);
	not #0 inv_14(RetC, net_16);
	not #0 inv_15(RetU, net_19);
	not #0 inv_16(CallC, net_11);
	not #0 inv_17(CallU, net_18);
	not #0 inv_18(BC, net_2);
	not #0 inv_19(BU, net_12);
	assign #0 net_12 = !(net_4 && net_17 && net_9 && enable);
	assign #0 net_6 = !(s[0] && s[1] && s[2] && enable);
	assign #0 net_20 = !(s[0] && s[1] && net_10 && enable);
	assign #0 net_16 = !(s[0] && net_14 && s[2] && enable);
	assign #0 net_19 = !(s[0] && net_5 && net_8 && enable);
	assign #0 net_11 = !(net_13 && s[1] && s[2] && enable);
	assign #0 net_18 = !(net_1 && s[1] && net_3 && enable);
	assign #0 net_2 = !(net_15 && net_7 && s[2] && enable);

endmodule		// BranchDecoder

module BranchEnable (BC, BE, BU, IR, N, P, T3, Z);
	input		BC;
	input		BU;
	input		N;
	input		P;
	input		T3;
	input		Z;
	input	[2:0]	IR;
	output		BE;
 
	wire		net_1;
	wire		net_2;
	wire		net_3;
	wire		net_4;
	wire		net_5;
	wire		net_6;
	wire		net_7;
	wire		net_8;
	wire		net_9;
 
	assign #0 net_5 = !(net_3 && BC);
	not #0 inv(net_8, net_5);
	not #0 inv_1(net_9, net_7);
	assign net_7 = !(net_8 || BU);
	assign #0 net_4 = !(net_9 && T3);
	assign #0 net_2 = !(IR[0] && Z);
	assign #0 net_6 = !(IR[1] && N);
	assign #0 net_1 = !(IR[2] && P);
	assign net_3 = !(net_2 || net_6 || net_1);
	not #0 inv_2(BE, net_4);

endmodule		// BranchEnable

module CallEnable (CE, CallC, CallU, IR, N, P, T3, Z);
	input		CallC;
	input		CallU;
	input		N;
	input		P;
	input		T3;
	input		Z;
	input	[2:0]	IR;
	output		CE;
 
	wire		net_1;
	wire		net_2;
	wire		net_3;
	wire		net_4;
	wire		net_5;
	wire		net_6;
	wire		net_7;
	wire		net_8;
	wire		net_9;
 
	assign #0 net_8 = !(net_9 && CallC);
	not #0 inv(net_5, net_8);
	not #0 inv_1(net_6, net_4);
	assign net_4 = !(net_5 || CallU);
	assign #0 net_7 = !(net_6 && T3);
	assign #0 net_2 = !(IR[0] && Z);
	assign #0 net_1 = !(IR[1] && N);
	assign #0 net_3 = !(IR[2] && P);
	assign net_9 = !(net_2 || net_1 || net_3);
	not #0 inv_2(CE, net_7);

endmodule		// CallEnable

module ReturnEnable (IR, N, P, RE, RetC, RetU, T3, Z);
	input		N;
	input		P;
	input		RetC;
	input		RetU;
	input		T3;
	input		Z;
	input	[2:0]	IR;
	output		RE;
 
	wire		net_1;
	wire		net_2;
	wire		net_3;
	wire		net_4;
	wire		net_5;
	wire		net_6;
	wire		net_7;
	wire		net_8;
	wire		net_9;
 
	assign #0 net_8 = !(net_9 && RetC);
	not #0 inv(net_5, net_8);
	not #0 inv_1(net_6, net_4);
	assign net_4 = !(net_5 || RetU);
	assign #0 net_7 = !(net_6 && T3);
	assign #0 net_2 = !(IR[0] && Z);
	assign #0 net_1 = !(IR[1] && N);
	assign #0 net_3 = !(IR[2] && P);
	assign net_9 = !(net_2 || net_1 || net_3);
	not #0 inv_2(RE, net_7);

endmodule		// ReturnEnable

module xor (in1, in2, out);
	input		in1;
	input		in2;
	output		out;
 
	wire		net_2;
	wire		net_3;
	wire		net_1;
 
	not #0 inv(net_1, in1);
	not #0 inv_1(out, net_2);
	not #0 inv_2(net_3, in2);
	xgate xgate(.in_L(net_1), .t2(net_2), .in(in1), .t1(in2));
	xgate xgate_1(.in(net_1), .t2(net_2), .t1(net_3), .in_L(in1));

endmodule		// xor

module Subtractor (A, Bin, Bout, D, F);
	input		A;
	input		Bin;
	input		F;
	output		Bout;
	output		D;
 
	wire		net_6;
	wire		net_2;
	wire		net_3;
	wire		net_4;
	wire		net_5;
	wire		net_1;
 
	xor xor(.out(net_6), .in2(A), .in1(F));
	xor xor_1(.in2(net_6), .out(D), .in1(Bin));
	assign #0 net_4 = !(Bin && F);
	assign #0 net_3 = !(Bin && net_2);
	assign #0 net_1 = !(F && net_5);
	assign Bout = !(net_4 || net_3 || net_1);
	not #0 inv(net_2, A);
	not #0 inv_1(net_5, A);

endmodule		// Subtractor

module Subtractor32bit (A, out, overflow);
	input	[31:0]	A;
	output		overflow;
	output	[31:0]	out;
 
	wire		net_28;
	wire		net_11;
	wire		net_30;
	wire		net_29;
	wire		net_12;
	wire		net_31;
	wire		net_13;
	wire		net_14;
	wire		net_15;
	wire		net_16;
	wire		net_17;
	wire		net_18;
	wire		net_1;
	wire		net_20;
	wire		net_19;
	wire		net_2;
	wire		net_21;
	wire		net_3;
	wire		net_22;
	wire		net_4;
	wire		net_23;
	wire		net_5;
	wire		net_24;
	wire		net_6;
	wire		net_25;
	wire		net_7;
	wire		net_26;
	wire		net_8;
	wire		net_27;
	wire		net_10;
	wire		net_9;
 
	Subtractor Subtractor(.Bout(net_3), .D(out[0]), .A(A[0]), .Bin(1'b0), 
		.F(1'b0));
	Subtractor Subtractor_1(.Bin(net_3), .Bout(net_30), .D(out[1]), 
		.A(A[1]), .F(1'b0));
	Subtractor Subtractor_2(.Bout(net_28), .Bin(net_30), .D(out[2]), 
		.A(A[2]), .F(1'b1));
	Subtractor Subtractor_3(.Bout(net_12), .Bin(net_28), .D(out[3]), 
		.A(A[3]), .F(1'b0));
	Subtractor Subtractor_4(.Bin(net_12), .Bout(net_18), .D(out[4]), 
		.A(A[4]), .F(1'b0));
	Subtractor Subtractor_5(.Bin(net_18), .Bout(net_19), .D(out[5]), 
		.A(A[5]), .F(1'b0));
	Subtractor Subtractor_6(.Bin(net_19), .Bout(net_27), .D(out[6]), 
		.A(A[6]), .F(1'b0));
	Subtractor Subtractor_7(.Bout(net_16), .Bin(net_27), .D(out[7]), 
		.A(A[7]), .F(1'b0));
	Subtractor Subtractor_8(.Bout(net_2), .Bin(net_16), .D(out[8]), 
		.A(A[8]), .F(1'b0));
	Subtractor Subtractor_9(.Bin(net_2), .Bout(net_4), .D(out[9]), 
		.A(A[9]), .F(1'b0));
	Subtractor Subtractor_10(.Bin(net_4), .Bout(net_9), .D(out[10]), 
		.A(A[10]), .F(1'b0));
	Subtractor Subtractor_11(.Bin(net_9), .Bout(net_22), .D(out[11]), 
		.A(A[11]), .F(1'b0));
	Subtractor Subtractor_12(.Bout(net_13), .Bin(net_22), .D(out[12]), 
		.A(A[12]), .F(1'b0));
	Subtractor Subtractor_13(.Bin(net_13), .Bout(net_15), .D(out[13]), 
		.A(A[13]), .F(1'b0));
	Subtractor Subtractor_14(.Bin(net_15), .Bout(net_23), .D(out[14]), 
		.A(A[14]), .F(1'b0));
	Subtractor Subtractor_15(.Bin(net_23), .Bout(net_24), .D(out[15]), 
		.A(A[15]), .F(1'b0));
	Subtractor Subtractor_16(.Bout(net_6), .Bin(net_24), .D(out[16]), 
		.A(A[16]), .F(1'b0));
	Subtractor Subtractor_17(.Bin(net_6), .Bout(net_29), .D(out[17]), 
		.A(A[17]), .F(1'b0));
	Subtractor Subtractor_18(.Bout(net_20), .Bin(net_29), .D(out[18]), 
		.A(A[18]), .F(1'b0));
	Subtractor Subtractor_19(.Bout(net_7), .Bin(net_20), .D(out[19]), 
		.A(A[19]), .F(1'b0));
	Subtractor Subtractor_20(.Bin(net_7), .Bout(net_14), .D(out[20]), 
		.A(A[20]), .F(1'b0));
	Subtractor Subtractor_21(.Bin(net_14), .Bout(net_21), .D(out[21]), 
		.A(A[21]), .F(1'b0));
	Subtractor Subtractor_22(.Bout(net_17), .Bin(net_21), .D(out[22]), 
		.A(A[22]), .F(1'b0));
	Subtractor Subtractor_23(.Bout(net_1), .Bin(net_17), .D(out[23]), 
		.A(A[23]), .F(1'b0));
	Subtractor Subtractor_24(.Bin(net_1), .Bout(net_25), .D(out[24]), 
		.A(A[24]), .F(1'b0));
	Subtractor Subtractor_25(.Bin(net_25), .Bout(net_26), .D(out[25]), 
		.A(A[25]), .F(1'b0));
	Subtractor Subtractor_26(.Bin(net_26), .Bout(net_31), .D(out[26]), 
		.A(A[26]), .F(1'b0));
	Subtractor Subtractor_27(.Bout(net_10), .Bin(net_31), .D(out[27]), 
		.A(A[27]), .F(1'b0));
	Subtractor Subtractor_28(.Bout(net_5), .Bin(net_10), .D(out[28]), 
		.A(A[28]), .F(1'b0));
	Subtractor Subtractor_29(.Bin(net_5), .Bout(net_8), .D(out[29]), 
		.A(A[29]), .F(1'b0));
	Subtractor Subtractor_30(.Bin(net_8), .Bout(net_11), .D(out[30]), 
		.A(A[30]), .F(1'b0));
	Subtractor Subtractor_31(.Bin(net_11), .D(out[31]), .A(A[31]), 
		.F(1'b0), .Bout(overflow));

endmodule		// Subtractor32bit

module BranchModule (BE, BRANCH_ENABLE, BRANCH_TARGET_ADDRESS, 
		BRANCH_TYPE, CE, IR, LS_ADDRESS, MDR_IN, N, P, R31_ADDRESS, RE, 
		SC_RESET_ENABLE, T3, T4, T6, Z, overflow);
	input		BRANCH_ENABLE;
	input		N;
	input		P;
	input		T3;
	input		T4;
	input		T6;
	input		Z;
	input	[2:0]	BRANCH_TYPE;
	input	[2:0]	IR;
	input	[31:0]	LS_ADDRESS;
	input	[31:0]	MDR_IN;
	input	[31:0]	R31_ADDRESS;
	output		BE;
	output		CE;
	output		RE;
	output		SC_RESET_ENABLE;
	output		overflow;
	output	[31:0]	BRANCH_TARGET_ADDRESS;
 
	wire		net_11;
	wire		net_12;
	wire		CE_int;
	wire	[1:0]	s;
	wire		net_1;
	wire		net_2;
	wire		net_3;
	wire		T3_int;
	wire		BE_int;
	wire		RE_int;
	wire		net_4;
	wire		net_5;
	wire	[31:0]	net_6;
	wire	[31:0]	latch;
	wire		net_7;
	wire		net_8;
	wire		net_10;
	wire		net_9;
 
	BranchDecoder BranchDecoder(.CallU(net_1), .BC(net_2), .CallC(net_4), 
		.BU(net_5), .RetU(net_10), .RetC(net_11), .enable(BRANCH_ENABLE), 
		.s(BRANCH_TYPE[2:0]));
	assign SC_RESET_ENABLE = !(BE_int || CE_int || RE_int);
	BranchEnable BranchEnable(.BC(net_2), .BU(net_5), .P(P), 
		.IR(IR[2:0]), .T3(1'b1), .BE(BE_int), .Z(Z), .N(N));
	CallEnable CallEnable(.CallU(net_1), .CallC(net_4), .P(P), 
		.CE(CE_int), .IR(IR[2:0]), .T3(1'b1), .Z(Z), .N(N));
	ReturnEnable ReturnEnable(.RetU(net_10), .RetC(net_11), .P(P), 
		.IR(IR[2:0]), .T3(1'b1), .RE(RE_int), .Z(Z), .N(N));
	Subtractor32bit Subtractor32bit(.out(net_6[31:0]), 
		.A(R31_ADDRESS[31:0]), .overflow(overflow));
	assign #0 net_12 = !(T3_int && RE_int);
	not #0 inv(net_7, net_12);
	DoubleInverter DoubleInverter(.out(RE), .in(RE_int));
	cell32trans cell32trans(.in(net_6[31:0]), .w(net_7), 
		.out(latch[31:0]));
	mux42132bbits mux42132bbits(.y(BRANCH_TARGET_ADDRESS[31:0]), 
		.s(s[1:0]), .b(R31_ADDRESS[31:0]), .a(LS_ADDRESS[31:0]), 
		.d(MDR_IN[31:0]), .c(latch[31:0]));
	DoubleInverter DoubleInverter_1(.out(CE), .in(CE_int));
	DoubleInverter DoubleInverter_2(.out(BE), .in(BE_int));
	assign #0 net_8 = !(CE_int && T3_int);
	assign #0 net_9 = !(RE_int && T4);
	assign #0 net_3 = !(RE_int && T6);
	assign s[0] = !(net_8 || net_3);
	assign s[1] = !(net_3 || net_9);
	DoubleInverter DoubleInverter_3(.in(T3), .out(T3_int));

endmodule		// BranchModule

module Mux5bit2to1 (a, b, s, y);
	input		s;
	input	[4:0]	a;
	input	[4:0]	b;
	output	[4:0]	y;
 
	wire		net_2;
	wire		net_1;
 
	Mux Mux(.s(net_1), .y(y[0]), .a(a[0]), .b(b[0]));
	Mux Mux_1(.s(net_1), .y(y[1]), .a(a[1]), .b(b[1]));
	Mux Mux_2(.s(net_1), .y(y[2]), .a(a[2]), .b(b[2]));
	Mux Mux_3(.s(net_1), .y(y[3]), .a(a[3]), .b(b[3]));
	not #0 inv(net_1, net_2);
	not #0 inv_1(net_2, s);
	Mux Mux_4(.s(net_1), .y(y[4]), .a(a[4]), .b(b[4]));

endmodule		// Mux5bit2to1

module Mux4to15bits (a, b, c, d, out, s);
	input	[4:0]	a;
	input	[4:0]	b;
	input	[4:0]	c;
	input	[4:0]	d;
	input	[1:0]	s;
	output	[4:0]	out;
 
	wire	[4:0]	net_2;
	wire	[4:0]	net_1;
 
	Mux5bit2to1 Mux5bit2to1(.y(net_1[4:0]), .a(a[4:0]), .b(b[4:0]), 
		.s(s[0]));
	Mux5bit2to1 Mux5bit2to1_1(.y(net_2[4:0]), .b(d[4:0]), .a(c[4:0]), 
		.s(s[0]));
	Mux5bit2to1 Mux5bit2to1_2(.a(net_1[4:0]), .b(net_2[4:0]), 
		.y(out[4:0]), .s(s[1]));

endmodule		// Mux4to15bits

module Mux5bits8to1 (a, b, c, d, e, f, g, h, out, s);
	input	[4:0]	a;
	input	[4:0]	b;
	input	[4:0]	c;
	input	[4:0]	d;
	input	[4:0]	e;
	input	[4:0]	f;
	input	[4:0]	g;
	input	[4:0]	h;
	input	[2:0]	s;
	output	[4:0]	out;
 
	wire	[4:0]	net_1;
	wire	[4:0]	net_2;
 
	Mux5bit2to1 Mux5bit2to1(.b(net_1[4:0]), .a(net_2[4:0]), .y(out[4:0]), 
		.s(s[2]));
	Mux4to15bits Mux4to15bits(.out(net_2[4:0]), .a(a[4:0]), .b(b[4:0]), 
		.s(s[1:0]), .c(c[4:0]), .d(d[4:0]));
	Mux4to15bits Mux4to15bits_1(.out(net_1[4:0]), .s(s[1:0]), .a(e[4:0]), 
		.b(f[4:0]), .c(g[4:0]), .d(h[4:0]));

endmodule		// Mux5bits8to1

module FinalProcessor (ALU_OVERFLOW, BRANCH_MODULE_OVERFLOW, CLOCK_IN, 
		LS_OVERFLOW, MAR_OUT, MDR_FROM_MEMORY, MDR_WE_FROM_MEMORY, 
		MDW_TO_MEMORY, MEMORY_READ, MEMORY_WRITE, PC_OVERFLOW, 
		STACKPOINTER_OVERFLOW);
	input		CLOCK_IN;
	input		MDR_WE_FROM_MEMORY;
	input	[31:0]	MDR_FROM_MEMORY;
	output		ALU_OVERFLOW;
	output		BRANCH_MODULE_OVERFLOW;
	output		LS_OVERFLOW;
	output		MEMORY_READ;
	output		MEMORY_WRITE;
	output		PC_OVERFLOW;
	output		STACKPOINTER_OVERFLOW;
	output	[31:0]	MAR_OUT;
	output	[31:0]	MDW_TO_MEMORY;
 
	wire		net_28;
	wire		net_30;
	wire		net_29;
	wire		net_31;
	wire	[1:0]	MDW_S;
	wire		net_32;
	wire		net_33;
	wire		net_34;
	wire		net_35;
	wire		net_36;
	wire	[31:0]	net_1;
	wire		net_37;
	wire		net_2;
	wire		net_38;
	wire		net_3;
	wire		net_40;
	wire	[4:0]	net_39;
	wire	[31:0]	MDR_OUT;
	wire	[31:0]	PC_OUT;
	wire	[4:0]	net_4;
	wire		net_41;
	wire		net_5;
	wire		net_6;
	wire		net_7;
	wire		net_8;
	wire		net_9;
	wire		BRANCH_UNIT_ACTIVATOR;
	wire	[7:0]	T;
	wire	[31:0]	LS_ADDRESS;
	wire	[31:0]	reg_out1;
	wire	[31:0]	reg_out2;
	wire		BE;
	wire		STORE_UNIT_ACTIVATOR;
	wire	[31:0]	IR_OUT;
	wire		CE;
	wire	[1:0]	ADDRESS_SOURCE_SELECT;
	wire		N_OUT;
	wire		P_OUT;
	wire		RE;
	wire		LOAD_UNIT_ACTIVATOR;
	wire	[2:0]	REG_FILE_S;
	wire		net_10;
	wire	[31:0]	net_11;
	wire		net_12;
	wire		Z_OUT;
	wire	[31:0]	BRANCH_TARGET_ADDRESS;
	wire		net_13;
	wire	[31:0]	net_14;
	wire		net_15;
	wire	[4:0]	net_16;
	wire		ALU_UNIT_ACTIVATOR;
	wire		net_17;
	wire	[4:0]	net_18;
	wire		net_20;
	wire		net_19;
	wire	[31:0]	ALU_RESULT;
	wire		net_21;
	wire		net_22;
	wire		net_23;
	wire	[1:0]	REG_WRITEADD_S;
	wire		net_24;
	wire		BRANCH_UNIT_RESET_SC;
	wire		net_25;
	wire		net_26;
	wire		net_27;
 
	DoubleInverter DoubleInverter(.in(net_27), .out(MEMORY_READ));
	assign #0 net_17 = !(ALU_UNIT_ACTIVATOR && IR_OUT[11] && T[4]);
	not #0 inv(net_6, net_17);
	ALU_UNIT ALU_UNIT(.PNZ_WE(net_6), .LATCH_WE(net_7), 
		.R1(reg_out1[31:0]), .R2(reg_out2[31:0]), .ALU_OP(IR_OUT[29:27]), 
		.N_OUT(N_OUT), .P_OUT(P_OUT), .ALU_OVERFLOW(ALU_OVERFLOW), 
		.Z_OUT(Z_OUT), .ALU_RESULT(ALU_RESULT[31:0]));
	assign #0 net_37 = !(T[4] && LOAD_UNIT_ACTIVATOR);
	DoubleInverter DoubleInverter_1(.in(net_25), .out(net_35));
	assign #0 net_25 = !(T[5] && STORE_UNIT_ACTIVATOR);
	assign #0 MDW_S[1] = !(T[4] && STORE_UNIT_ACTIVATOR);
	assign #0 net_7 = !(T[3] && ALU_UNIT_ACTIVATOR);
	LoadStoreModule LoadStoreModule(.LS_OVERFLOW(LS_OVERFLOW), .T0(T[0]), 
		.T3(T[3]), .LS_ADDRESS(LS_ADDRESS[31:0]), 
		.R_BASE_VALUE(reg_out2[31:0]), .STORE(STORE_UNIT_ACTIVATOR), 
		.OFFSET(IR_OUT[16:0]), .S(ADDRESS_SOURCE_SELECT[1:0]), 
		.LOAD(LOAD_UNIT_ACTIVATOR));
	assign #0 net_28 = !(BE && T[3]);
	assign #0 net_2 = !(LOAD_UNIT_ACTIVATOR && T[3]);
	assign #0 net_32 = !(STORE_UNIT_ACTIVATOR && T[3]);
	assign #0 net_13 = !(CE && T[3]);
	assign #0 net_21 = !(CE && T[5]);
	assign #0 net_12 = !(RE && T[4]);
	assign #0 net_23 = !(RE && T[6]);
	assign net_41 = !(net_2 || net_32 || net_28 || net_13 || net_21 || 
		net_12 || net_23);
	assign net_8 = !(net_28 || net_13 || net_21 || net_12 || net_23);
	controlunit controlunit(.MDW_WE(net_3), .SC_RESET(net_5), 
		.BRANCH_ENABLE(net_8), .MDW_IN(net_14[31:0]), .MAR_WE(net_41), 
		.CLOCK(CLOCK_IN), .MDW_OUT(MDW_TO_MEMORY[31:0]), 
		.MDR_OUT(MDR_OUT[31:0]), .PC_OUT(PC_OUT[31:0]), 
		.MAR_OUT(MAR_OUT[31:0]), 
		.BRANCH_UNIT_ACTIVATOR(BRANCH_UNIT_ACTIVATOR), .T_OUT(T[7:0]), 
		.STORE_UNIT_ADDRESS(LS_ADDRESS[31:0]), 
		.LOAD_UNIT_ADDRESS(LS_ADDRESS[31:0]), 
		.STORE_UNIT_ACTIVATOR(STORE_UNIT_ACTIVATOR), .IR_OUT(IR_OUT[31:0]), 
		.MDR_IN(MDR_FROM_MEMORY[31:0]), 
		.ADDRESS_SOURCE_SELECT(ADDRESS_SOURCE_SELECT[1:0]), 
		.MDR_WE(MDR_WE_FROM_MEMORY), 
		.LOAD_UNIT_ACTIVATOR(LOAD_UNIT_ACTIVATOR), 
		.BRANCH_TARGET(BRANCH_TARGET_ADDRESS[31:0]), 
		.ALU_UNIT_ACTIVATOR(ALU_UNIT_ACTIVATOR), .PC_OVERFLOW(PC_OVERFLOW));
	assign #0 MDW_S[0] = !(T[4] && CE);
	assign net_3 = !(MDW_S[1] || MDW_S[0]);
	mux42132bbits mux42132bbits(.y(net_14[31:0]), 
		.a({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), 
		.d({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), 
		.s(MDW_S[1:0]), .c(PC_OUT[31:0]), .b(reg_out1[31:0]));
	DoubleInverter DoubleInverter_2(.out(net_36), .in(net_38));
	assign #0 net_38 = !(T[5] && CE);
	assign MEMORY_WRITE = !(net_35 || net_36);
	assign net_27 = !(net_26 || net_20 || net_37);
	assign #0 net_20 = !(T[5] && CE);
	not #0 inv_1(net_26, T[1]);
	Register_file_32bits Register_file_32bits(.data(net_1[31:0]), 
		.address_read1(net_4[4:0]), .address_write(net_16[4:0]), 
		.write_enable(net_30), .OUT1(reg_out1[31:0]), .OUT2(reg_out2[31:0]), 
		.address_read2(IR_OUT[21:17]));
	assign #0 net_34 = !(T[4] && ALU_UNIT_ACTIVATOR);
	assign #0 net_33 = !(T[5] && LOAD_UNIT_ACTIVATOR);
	assign #0 net_31 = !(T[4] && CE);
	assign net_30 = !(net_34 || net_33 || net_31);
	assign #0 net_15 = !(T[5] && ALU_UNIT_ACTIVATOR);
	assign #0 net_29 = !(T[6] && LOAD_UNIT_ACTIVATOR);
	assign #0 net_10 = !(T[6] && STORE_UNIT_ACTIVATOR);
	assign #0 net_19 = !(T[4] && BE);
	assign #0 net_24 = !(T[6] && CE);
	assign #0 net_22 = !(T[7] && RE);
	assign net_5 = !(BRANCH_UNIT_RESET_SC || net_22 || net_24 || net_19 
		|| net_10 || net_29 || net_15);
	FiveOnes FiveOnes(.out(net_39[4:0]));
	assign net_40 = !(LOAD_UNIT_ACTIVATOR || STORE_UNIT_ACTIVATOR);
	not #0 inv_2(REG_FILE_S[1], net_40);
	DoubleInverter DoubleInverter_3(.out(REG_FILE_S[0]), 
		.in(ALU_UNIT_ACTIVATOR));
	DoubleInverter DoubleInverter_4(.in(BRANCH_UNIT_ACTIVATOR), 
		.out(REG_FILE_S[2]));
	Mux32Bit8to1 Mux32Bit8to1(.out(net_1[31:0]), .E(net_11[31:0]), 
		.D({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), 
		.F({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), 
		.G({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), 
		.H({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), 
		.A({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), 
		.C(MDR_OUT[31:0]), .s(REG_FILE_S[2:0]), .B(ALU_RESULT[31:0]));
	FiveOnes FiveOnes_1(.out(net_18[4:0]));
	pcincrement pcincrement(.s(net_11[31:0]), 
		.overflow(STACKPOINTER_OVERFLOW), .a(MAR_OUT[31:0]));
	BranchModule BranchModule(.MDR_IN(MDR_OUT[31:0]), 
		.BRANCH_ENABLE(BRANCH_UNIT_ACTIVATOR), .T3(T[3]), .T6(T[6]), 
		.T4(T[4]), .LS_ADDRESS(LS_ADDRESS[31:0]), 
		.R31_ADDRESS(reg_out1[31:0]), .BE(BE), .IR(IR_OUT[24:22]), 
		.BRANCH_TYPE(IR_OUT[28:26]), .CE(CE), .N(N_OUT), .P(P_OUT), .RE(RE), 
		.overflow(BRANCH_MODULE_OVERFLOW), .Z(Z_OUT), 
		.BRANCH_TARGET_ADDRESS(BRANCH_TARGET_ADDRESS[31:0]), 
		.SC_RESET_ENABLE(BRANCH_UNIT_RESET_SC));
	Mux4to15bits Mux4to15bits(.out(net_16[4:0]), .c(net_18[4:0]), 
		.a({1'b0,1'b0,1'b0,1'b0,1'b0}), .d({1'b0,1'b0,1'b0,1'b0,1'b0}), 
		.b(IR_OUT[26:22]), .s(REG_WRITEADD_S[1:0]));
	not #0 inv_3(REG_WRITEADD_S[0], net_9);
	assign net_9 = !(LOAD_UNIT_ACTIVATOR || STORE_UNIT_ACTIVATOR || 
		ALU_UNIT_ACTIVATOR);
	DoubleInverter DoubleInverter_5(.in(BRANCH_UNIT_ACTIVATOR), 
		.out(REG_WRITEADD_S[1]));
	Mux5bits8to1 Mux5bits8to1(.out(net_4[4:0]), .e(net_39[4:0]), 
		.a({1'b0,1'b0,1'b0,1'b0,1'b0}), .d({1'b0,1'b0,1'b0,1'b0,1'b0}), 
		.f({1'b0,1'b0,1'b0,1'b0,1'b0}), .g({1'b0,1'b0,1'b0,1'b0,1'b0}), 
		.h({1'b0,1'b0,1'b0,1'b0,1'b0}), .b(IR_OUT[16:12]), 
		.c(IR_OUT[26:22]), .s(REG_FILE_S[2:0]));
	Inverters32Bit Inverters32Bit(.in(MAR_OUT[31:0]), 
		.out(MAR_OUT[31:0]));

endmodule		// FinalProcessor

